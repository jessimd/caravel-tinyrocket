module SRAM1RW4096x8 (
	A,
	CE,
	I,
	O,
	CSB,
	OEB,
	WEB
);
	input [11:0] A;
	input CE;
	input [7:0] I;
	output wire [7:0] O;
	input CSB;
	input OEB;
	input WEB;
	wire [10:0] addr0;
	wire [3:0] wmask0;
	wire [32:0] din0;
	wire [32:0] dout0;
	wire [1:0] index;
	assign index = A[1:0];
	assign din0[index * 8+:8] = I;
	assign O = dout0[index * 8+:8];
	assign addr0 = {1'b0, A[11:2]};
	assign wmask0 = {{index[1] && !index[0]}, {index[1] && index[0]}, {!index[1] && index[0]}, {!index[1] && !index[0]}};
	wire vccd1;
	wire vssd1;
	sky130_sram_4kbyte_1rw_32x1024_8 sram_4096x8(
		.vccd1(vccd1),
		.vssd1(vssd1),
		.clk0(CE),
		.csb0(CSB),
		.web0(WEB),
		.wmask0(wmask0),
		.addr0(addr0),
		.din0(din0),
		.dout0(dout0)
	);
endmodule
module SRAM1RW64x21 (
	A,
	CE,
	I,
	O,
	CSB,
	OEB,
	WEB
);
	input [5:0] A;
	input CE;
	input [20:0] I;
	output wire [20:0] O;
	input CSB;
	input OEB;
	input WEB;
	wire vccd1;
	wire vssd1;
	sky130_sram_0kbytes_1rw_21x64_21 sram_64x21(
		.vccd1(vccd1),
		.vssd1(vssd1),
		.clk0(CE),
		.csb0(CSB),
		.web0(WEB),
		.addr0(A),
		.din0(I),
		.dout0(O)
	);
endmodule
module SRAM1RW1024x32 (
	A,
	CE,
	I,
	O,
	CSB,
	OEB,
	WEB
);
	input [9:0] A;
	input CE;
	input [31:0] I;
	output wire [31:0] O;
	input CSB;
	input OEB;
	input WEB;
	wire vccd1;
	wire vssd1;
	sky130_sram_4kbytes_1rw_32x1024_32 sram_1024x32(
		.vccd1(vccd1),
		.vssd1(vssd1),
		.clk0(CE),
		.csb0(CSB),
		.web0(WEB),
		.addr0(A),
		.din0(I),
		.dout0(O)
	);
endmodule
module SRAM1RW1024x37 (
	A,
	CE,
	I,
	O,
	CSB,
	OEB,
	WEB
);
	input [9:0] A;
	input CE;
	input [36:0] I;
	output wire [36:0] O;
	input CSB;
	input OEB;
	input WEB;
	wire vccd1;
	wire vssd1;
	sky130_sram_5kbytes_1rw_37x1024_37 sram_1024x37(
		.vccd1(vccd1),
		.vssd1(vssd1),
		.clk0(CE),
		.csb0(CSB),
		.web0(WEB),
		.addr0(A),
		.din0(I),
		.dout0(O)
	);
endmodule
module sky130_sram_4kbytes_1rw_32x1024_32 (
	vccd1,
	vssd1,
	clk0,
	csb0,
	web0,
	spare_wen0,
	addr0,
	din0,
	dout0
);
	inout vccd1;
	inout vssd1;
	input clk0;
	input csb0;
	input web0;
	input [10:0] addr0;
	input spare_wen0;
	input [32:0] din0;
	output wire [32:0] dout0;
endmodule
module data_arrays_0_ext (
	RW0_addr,
	RW0_clk,
	RW0_wdata,
	RW0_rdata,
	RW0_en,
	RW0_wmode,
	RW0_wmask
);
	input [11:0] RW0_addr;
	input RW0_clk;
	input [31:0] RW0_wdata;
	output wire [31:0] RW0_rdata;
	input RW0_en;
	input RW0_wmode;
	input [3:0] RW0_wmask;
	wire [11:0] mem_0_0_A;
	wire mem_0_0_CE;
	wire [7:0] mem_0_0_I;
	wire [7:0] mem_0_0_O;
	wire mem_0_0_CSB;
	wire mem_0_0_OEB;
	wire mem_0_0_WEB;
	wire [11:0] mem_0_1_A;
	wire mem_0_1_CE;
	wire [7:0] mem_0_1_I;
	wire [7:0] mem_0_1_O;
	wire mem_0_1_CSB;
	wire mem_0_1_OEB;
	wire mem_0_1_WEB;
	wire [11:0] mem_0_2_A;
	wire mem_0_2_CE;
	wire [7:0] mem_0_2_I;
	wire [7:0] mem_0_2_O;
	wire mem_0_2_CSB;
	wire mem_0_2_OEB;
	wire mem_0_2_WEB;
	wire [11:0] mem_0_3_A;
	wire mem_0_3_CE;
	wire [7:0] mem_0_3_I;
	wire [7:0] mem_0_3_O;
	wire mem_0_3_CSB;
	wire mem_0_3_OEB;
	wire mem_0_3_WEB;
	wire [7:0] RW0_rdata_0_0 = mem_0_0_O;
	wire [7:0] RW0_rdata_0_1 = mem_0_1_O;
	wire [7:0] RW0_rdata_0_2 = mem_0_2_O;
	wire [7:0] RW0_rdata_0_3 = mem_0_3_O;
	wire [15:0] _GEN_0 = {RW0_rdata_0_1, RW0_rdata_0_0};
	wire [23:0] _GEN_1 = {RW0_rdata_0_2, RW0_rdata_0_1, RW0_rdata_0_0};
	wire [31:0] RW0_rdata_0 = {RW0_rdata_0_3, RW0_rdata_0_2, RW0_rdata_0_1, RW0_rdata_0_0};
	wire [15:0] _GEN_2 = {RW0_rdata_0_1, RW0_rdata_0_0};
	wire [23:0] _GEN_3 = {RW0_rdata_0_2, RW0_rdata_0_1, RW0_rdata_0_0};
	wire _GEN_4 = ~RW0_wmode;
	wire _GEN_5 = ~RW0_wmode & RW0_en;
	wire _GEN_6 = RW0_wmask[0];
	wire _GEN_7 = RW0_wmode & RW0_wmask[0];
	wire _GEN_8 = ~RW0_wmode;
	wire _GEN_9 = ~RW0_wmode & RW0_en;
	wire _GEN_10 = RW0_wmask[1];
	wire _GEN_11 = RW0_wmode & RW0_wmask[1];
	wire _GEN_12 = ~RW0_wmode;
	wire _GEN_13 = ~RW0_wmode & RW0_en;
	wire _GEN_14 = RW0_wmask[2];
	wire _GEN_15 = RW0_wmode & RW0_wmask[2];
	wire _GEN_16 = ~RW0_wmode;
	wire _GEN_17 = ~RW0_wmode & RW0_en;
	wire _GEN_18 = RW0_wmask[3];
	wire _GEN_19 = RW0_wmode & RW0_wmask[3];
	SRAM1RW4096x8 mem_0_0(
		.A(mem_0_0_A),
		.CE(mem_0_0_CE),
		.I(mem_0_0_I),
		.O(mem_0_0_O),
		.CSB(mem_0_0_CSB),
		.OEB(mem_0_0_OEB),
		.WEB(mem_0_0_WEB)
	);
	SRAM1RW4096x8 mem_0_1(
		.A(mem_0_1_A),
		.CE(mem_0_1_CE),
		.I(mem_0_1_I),
		.O(mem_0_1_O),
		.CSB(mem_0_1_CSB),
		.OEB(mem_0_1_OEB),
		.WEB(mem_0_1_WEB)
	);
	SRAM1RW4096x8 mem_0_2(
		.A(mem_0_2_A),
		.CE(mem_0_2_CE),
		.I(mem_0_2_I),
		.O(mem_0_2_O),
		.CSB(mem_0_2_CSB),
		.OEB(mem_0_2_OEB),
		.WEB(mem_0_2_WEB)
	);
	SRAM1RW4096x8 mem_0_3(
		.A(mem_0_3_A),
		.CE(mem_0_3_CE),
		.I(mem_0_3_I),
		.O(mem_0_3_O),
		.CSB(mem_0_3_CSB),
		.OEB(mem_0_3_OEB),
		.WEB(mem_0_3_WEB)
	);
	assign RW0_rdata = {RW0_rdata_0_3, _GEN_1};
	assign mem_0_0_A = RW0_addr;
	assign mem_0_0_CE = RW0_clk;
	assign mem_0_0_I = RW0_wdata[7:0];
	assign mem_0_0_CSB = ~RW0_en;
	assign mem_0_0_OEB = ~(~RW0_wmode & RW0_en);
	assign mem_0_0_WEB = ~(RW0_wmode & RW0_wmask[0]);
	assign mem_0_1_A = RW0_addr;
	assign mem_0_1_CE = RW0_clk;
	assign mem_0_1_I = RW0_wdata[15:8];
	assign mem_0_1_CSB = ~RW0_en;
	assign mem_0_1_OEB = ~(~RW0_wmode & RW0_en);
	assign mem_0_1_WEB = ~(RW0_wmode & RW0_wmask[1]);
	assign mem_0_2_A = RW0_addr;
	assign mem_0_2_CE = RW0_clk;
	assign mem_0_2_I = RW0_wdata[23:16];
	assign mem_0_2_CSB = ~RW0_en;
	assign mem_0_2_OEB = ~(~RW0_wmode & RW0_en);
	assign mem_0_2_WEB = ~(RW0_wmode & RW0_wmask[2]);
	assign mem_0_3_A = RW0_addr;
	assign mem_0_3_CE = RW0_clk;
	assign mem_0_3_I = RW0_wdata[31:24];
	assign mem_0_3_CSB = ~RW0_en;
	assign mem_0_3_OEB = ~(~RW0_wmode & RW0_en);
	assign mem_0_3_WEB = ~(RW0_wmode & RW0_wmask[3]);
endmodule
module tag_array_ext (
	RW0_addr,
	RW0_clk,
	RW0_wdata,
	RW0_rdata,
	RW0_en,
	RW0_wmode,
	RW0_wmask
);
	input [5:0] RW0_addr;
	input RW0_clk;
	input [20:0] RW0_wdata;
	output wire [20:0] RW0_rdata;
	input RW0_en;
	input RW0_wmode;
	input RW0_wmask;
	wire [5:0] mem_0_0_A;
	wire mem_0_0_CE;
	wire [20:0] mem_0_0_I;
	wire [20:0] mem_0_0_O;
	wire mem_0_0_CSB;
	wire mem_0_0_OEB;
	wire mem_0_0_WEB;
	wire [20:0] RW0_rdata_0_0 = mem_0_0_O;
	wire [20:0] RW0_rdata_0 = RW0_rdata_0_0;
	wire _GEN_0 = ~RW0_wmode;
	wire _GEN_1 = ~RW0_wmode & RW0_en;
	wire _GEN_2 = RW0_wmode & RW0_wmask;
	SRAM1RW64x21 mem_0_0(
		.A(mem_0_0_A),
		.CE(mem_0_0_CE),
		.I(mem_0_0_I),
		.O(mem_0_0_O),
		.CSB(mem_0_0_CSB),
		.OEB(mem_0_0_OEB),
		.WEB(mem_0_0_WEB)
	);
	assign RW0_rdata = mem_0_0_O;
	assign mem_0_0_A = RW0_addr;
	assign mem_0_0_CE = RW0_clk;
	assign mem_0_0_I = RW0_wdata;
	assign mem_0_0_CSB = ~RW0_en;
	assign mem_0_0_OEB = ~(~RW0_wmode & RW0_en);
	assign mem_0_0_WEB = ~(RW0_wmode & RW0_wmask);
endmodule
module data_arrays_0_0_ext (
	RW0_addr,
	RW0_clk,
	RW0_wdata,
	RW0_rdata,
	RW0_en,
	RW0_wmode,
	RW0_wmask
);
	input [9:0] RW0_addr;
	input RW0_clk;
	input [31:0] RW0_wdata;
	output wire [31:0] RW0_rdata;
	input RW0_en;
	input RW0_wmode;
	input RW0_wmask;
	wire [9:0] mem_0_0_A;
	wire mem_0_0_CE;
	wire [31:0] mem_0_0_I;
	wire [31:0] mem_0_0_O;
	wire mem_0_0_CSB;
	wire mem_0_0_OEB;
	wire mem_0_0_WEB;
	wire [31:0] RW0_rdata_0_0 = mem_0_0_O;
	wire [31:0] RW0_rdata_0 = RW0_rdata_0_0;
	wire _GEN_0 = ~RW0_wmode;
	wire _GEN_1 = ~RW0_wmode & RW0_en;
	wire _GEN_2 = RW0_wmode & RW0_wmask;
	SRAM1RW1024x32 mem_0_0(
		.A(mem_0_0_A),
		.CE(mem_0_0_CE),
		.I(mem_0_0_I),
		.O(mem_0_0_O),
		.CSB(mem_0_0_CSB),
		.OEB(mem_0_0_OEB),
		.WEB(mem_0_0_WEB)
	);
	assign RW0_rdata = mem_0_0_O;
	assign mem_0_0_A = RW0_addr;
	assign mem_0_0_CE = RW0_clk;
	assign mem_0_0_I = RW0_wdata;
	assign mem_0_0_CSB = ~RW0_en;
	assign mem_0_0_OEB = ~(~RW0_wmode & RW0_en);
	assign mem_0_0_WEB = ~(RW0_wmode & RW0_wmask);
endmodule
module l2_tlb_ram_ext (
	RW0_addr,
	RW0_clk,
	RW0_wdata,
	RW0_rdata,
	RW0_en,
	RW0_wmode
);
	input [9:0] RW0_addr;
	input RW0_clk;
	input [36:0] RW0_wdata;
	output wire [36:0] RW0_rdata;
	input RW0_en;
	input RW0_wmode;
	wire [9:0] mem_0_0_A;
	wire mem_0_0_CE;
	wire [36:0] mem_0_0_I;
	wire [36:0] mem_0_0_O;
	wire mem_0_0_CSB;
	wire mem_0_0_OEB;
	wire mem_0_0_WEB;
	wire [36:0] RW0_rdata_0_0 = mem_0_0_O;
	wire [36:0] RW0_rdata_0 = RW0_rdata_0_0;
	wire _GEN_0 = ~RW0_wmode;
	wire _GEN_1 = ~RW0_wmode & RW0_en;
	SRAM1RW1024x37 mem_0_0(
		.A(mem_0_0_A),
		.CE(mem_0_0_CE),
		.I(mem_0_0_I),
		.O(mem_0_0_O),
		.CSB(mem_0_0_CSB),
		.OEB(mem_0_0_OEB),
		.WEB(mem_0_0_WEB)
	);
	assign RW0_rdata = mem_0_0_O;
	assign mem_0_0_A = RW0_addr;
	assign mem_0_0_CE = RW0_clk;
	assign mem_0_0_I = RW0_wdata;
	assign mem_0_0_CSB = ~RW0_en;
	assign mem_0_0_OEB = ~(~RW0_wmode & RW0_en);
	assign mem_0_0_WEB = ~RW0_wmode;
endmodule
module GenericAnalogIOCell (
	pad,
	core
);
	inout pad;
	inout core;
	assign core = 1'bz;
	assign pad = core;
endmodule
module GenericDigitalGPIOCell (
	pad,
	i,
	ie,
	o,
	oe
);
	inout pad;
	output wire i;
	input ie;
	input o;
	input oe;
	assign pad = (oe ? o : 1'bz);
	assign i = (ie ? pad : 1'b0);
endmodule
module GenericDigitalInIOCell (
	pad,
	i,
	ie
);
	input pad;
	output wire i;
	input ie;
	assign i = (ie ? pad : 1'b0);
endmodule
module GenericDigitalOutIOCell (
	pad,
	o,
	oe
);
	output wire pad;
	input o;
	input oe;
	assign pad = (oe ? o : 1'bz);
endmodule
module ClockDividerN (
	clk_out,
	clk_in
);
	parameter DIV = 1;
	output reg clk_out = 1'b0;
	input clk_in;
	localparam CWIDTH = $clog2(DIV);
	localparam LOW_CYCLES = DIV / 2;
	localparam HIGH_TRANSITION = LOW_CYCLES - 1;
	localparam LOW_TRANSITION = DIV - 1;
	generate
		if (DIV == 1) begin : genblk1
			always @(clk_in) clk_out = clk_in;
		end
		else begin : genblk1
			reg [CWIDTH - 1:0] count = HIGH_TRANSITION[CWIDTH - 1:0];
			always @(posedge clk_in)
				if (count == LOW_TRANSITION[CWIDTH - 1:0]) begin
					clk_out = 1'b0;
					count <= 1'sb0;
				end
				else begin
					if (count == HIGH_TRANSITION[CWIDTH - 1:0])
						clk_out = 1'b1;
					count <= count + 1'b1;
				end
		end
	endgenerate
endmodule
module plusarg_reader (out);
	parameter FORMAT = "borked=%d";
	parameter WIDTH = 1;
	parameter [WIDTH - 1:0] DEFAULT = 0;
	output wire [WIDTH - 1:0] out;
	assign out = DEFAULT;
endmodule
module EICG_wrapper (
	out,
	en,
	test_en,
	in
);
	output wire out;
	input en;
	input test_en;
	input in;
	reg en_latched;
	always @(*)
		if (!in)
			en_latched = en || test_en;
	assign out = en_latched && in;
endmodule
module sky130_sram_5kbytes_1rw_37x1024_37 (
	clk0,
	csb0,
	web0,
	spare_wen0,
	addr0,
	din0,
	dout0,
	vccd1,
	vssd1
);
	input clk0;
	input csb0;
	input web0;
	input [9:0] addr0;
	input spare_wen0;
	input [36:0] din0;
	output wire [36:0] dout0;
	inout vccd1;
	inout vssd1;
endmodule
module IntXbar (
	auto_int_in_0,
	auto_int_out_0
);
	input auto_int_in_0;
	output wire auto_int_out_0;
	assign auto_int_out_0 = auto_int_in_0;
endmodule
module InterruptBusWrapper (
	auto_int_bus_int_in_0,
	auto_int_bus_int_out_0
);
	input auto_int_bus_int_in_0;
	output wire auto_int_bus_int_out_0;
	wire int_bus_auto_int_in_0;
	wire int_bus_auto_int_out_0;
	IntXbar int_bus(
		.auto_int_in_0(int_bus_auto_int_in_0),
		.auto_int_out_0(int_bus_auto_int_out_0)
	);
	assign auto_int_bus_int_out_0 = int_bus_auto_int_out_0;
	assign int_bus_auto_int_in_0 = auto_int_bus_int_in_0;
endmodule
module ClockGroupAggregator (
	auto_in_member_subsystem_sbus_0_clock,
	auto_in_member_subsystem_sbus_0_reset,
	auto_out_member_subsystem_sbus_0_clock,
	auto_out_member_subsystem_sbus_0_reset
);
	input auto_in_member_subsystem_sbus_0_clock;
	input auto_in_member_subsystem_sbus_0_reset;
	output wire auto_out_member_subsystem_sbus_0_clock;
	output wire auto_out_member_subsystem_sbus_0_reset;
	assign auto_out_member_subsystem_sbus_0_clock = auto_in_member_subsystem_sbus_0_clock;
	assign auto_out_member_subsystem_sbus_0_reset = auto_in_member_subsystem_sbus_0_reset;
endmodule
module ClockGroup (
	auto_in_member_subsystem_sbus_0_clock,
	auto_in_member_subsystem_sbus_0_reset,
	auto_out_clock,
	auto_out_reset
);
	input auto_in_member_subsystem_sbus_0_clock;
	input auto_in_member_subsystem_sbus_0_reset;
	output wire auto_out_clock;
	output wire auto_out_reset;
	assign auto_out_clock = auto_in_member_subsystem_sbus_0_clock;
	assign auto_out_reset = auto_in_member_subsystem_sbus_0_reset;
endmodule
module FixedClockBroadcast (
	auto_in_clock,
	auto_in_reset,
	auto_out_2_clock,
	auto_out_2_reset,
	auto_out_0_clock,
	auto_out_0_reset
);
	input auto_in_clock;
	input auto_in_reset;
	output wire auto_out_2_clock;
	output wire auto_out_2_reset;
	output wire auto_out_0_clock;
	output wire auto_out_0_reset;
	assign auto_out_2_clock = auto_in_clock;
	assign auto_out_2_reset = auto_in_reset;
	assign auto_out_0_clock = auto_in_clock;
	assign auto_out_0_reset = auto_in_reset;
endmodule
module TLMonitor (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = ~io_in_a_bits_source;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_5 = ~_source_ok_T;
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_15 = io_in_a_bits_opcode == 3'h6;
	wire _T_17 = io_in_a_bits_size <= 4'hc;
	wire _T_20 = _T_17 & _source_ok_T;
	wire [32:0] _T_26 = $signed(_T_7) & -33'sh000005000;
	wire _T_27 = $signed(_T_26) == 33'sh000000000;
	wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_29 = {1'b0, $signed(_T_28)};
	wire [32:0] _T_31 = $signed(_T_29) & -33'sh000001000;
	wire _T_32 = $signed(_T_31) == 33'sh000000000;
	wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [32:0] _T_36 = $signed(_T_34) & -33'sh000010000;
	wire _T_37 = $signed(_T_36) == 33'sh000000000;
	wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_39 = {1'b0, $signed(_T_38)};
	wire [32:0] _T_41 = $signed(_T_39) & -33'sh000010000;
	wire _T_42 = $signed(_T_41) == 33'sh000000000;
	wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_44 = {1'b0, $signed(_T_43)};
	wire [32:0] _T_46 = $signed(_T_44) & -33'sh000011000;
	wire _T_47 = $signed(_T_46) == 33'sh000000000;
	wire [31:0] _T_48 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_49 = {1'b0, $signed(_T_48)};
	wire [32:0] _T_51 = $signed(_T_49) & -33'sh000010000;
	wire _T_52 = $signed(_T_51) == 33'sh000000000;
	wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_54 = {1'b0, $signed(_T_53)};
	wire [32:0] _T_56 = $signed(_T_54) & -33'sh004000000;
	wire _T_57 = $signed(_T_56) == 33'sh000000000;
	wire [31:0] _T_58 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_59 = {1'b0, $signed(_T_58)};
	wire [32:0] _T_61 = $signed(_T_59) & -33'sh000001000;
	wire _T_62 = $signed(_T_61) == 33'sh000000000;
	wire [31:0] _T_63 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_64 = {1'b0, $signed(_T_63)};
	wire [32:0] _T_66 = $signed(_T_64) & -33'sh000001000;
	wire _T_67 = $signed(_T_66) == 33'sh000000000;
	wire [31:0] _T_68 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_69 = {1'b0, $signed(_T_68)};
	wire [32:0] _T_71 = $signed(_T_69) & -33'sh000004000;
	wire _T_72 = $signed(_T_71) == 33'sh000000000;
	wire _T_167 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_171 = ~io_in_a_bits_mask;
	wire _T_172 = _T_171 == 4'h0;
	wire _T_176 = ~io_in_a_bits_corrupt;
	wire _T_180 = io_in_a_bits_opcode == 3'h7;
	wire _T_336 = io_in_a_bits_param != 3'h0;
	wire _T_349 = io_in_a_bits_opcode == 3'h4;
	wire _T_368 = _T_17 & _T_32;
	wire _T_370 = io_in_a_bits_size <= 4'h6;
	wire _T_425 = (((((((_T_27 | _T_37) | _T_42) | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_426 = _T_370 & _T_425;
	wire _T_428 = _T_368 | _T_426;
	wire _T_438 = io_in_a_bits_param == 3'h0;
	wire _T_442 = io_in_a_bits_mask == mask;
	wire _T_450 = io_in_a_bits_opcode == 3'h0;
	wire _T_511 = (((((_T_27 | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_512 = _T_370 & _T_511;
	wire _T_527 = _T_368 | _T_512;
	wire _T_529 = _T_20 & _T_527;
	wire _T_547 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_640 = ~mask;
	wire [3:0] _T_641 = io_in_a_bits_mask & _T_640;
	wire _T_642 = _T_641 == 4'h0;
	wire _T_646 = io_in_a_bits_opcode == 3'h2;
	wire _T_654 = io_in_a_bits_size <= 4'h2;
	wire _T_703 = ((((((_T_27 | _T_32) | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_704 = _T_654 & _T_703;
	wire _T_720 = _T_20 & _T_704;
	wire _T_730 = io_in_a_bits_param <= 3'h4;
	wire _T_738 = io_in_a_bits_opcode == 3'h3;
	wire _T_822 = io_in_a_bits_param <= 3'h3;
	wire _T_830 = io_in_a_bits_opcode == 3'h5;
	wire _T_904 = _T_20 & _T_368;
	wire _T_914 = io_in_a_bits_param <= 3'h1;
	wire _T_926 = io_in_d_bits_opcode <= 3'h6;
	wire _T_930 = io_in_d_bits_opcode == 3'h6;
	wire _T_934 = io_in_d_bits_size >= 4'h2;
	wire _T_938 = io_in_d_bits_param == 2'h0;
	wire _T_942 = ~io_in_d_bits_corrupt;
	wire _T_946 = ~io_in_d_bits_denied;
	wire _T_950 = io_in_d_bits_opcode == 3'h4;
	wire _T_961 = io_in_d_bits_param <= 2'h2;
	wire _T_965 = io_in_d_bits_param != 2'h2;
	wire _T_978 = io_in_d_bits_opcode == 3'h5;
	wire _T_998 = _T_946 | io_in_d_bits_corrupt;
	wire _T_1007 = io_in_d_bits_opcode == 3'h0;
	wire _T_1024 = io_in_d_bits_opcode == 3'h1;
	wire _T_1042 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg source;
	reg [31:0] address;
	wire _T_1072 = io_in_a_valid & ~a_first;
	wire _T_1073 = io_in_a_bits_opcode == opcode;
	wire _T_1077 = io_in_a_bits_param == param;
	wire _T_1081 = io_in_a_bits_size == size;
	wire _T_1085 = io_in_a_bits_source == source;
	wire _T_1089 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg sink;
	reg denied;
	wire _T_1096 = io_in_d_valid & ~d_first;
	wire _T_1097 = io_in_d_bits_opcode == opcode_1;
	wire _T_1101 = io_in_d_bits_param == param_1;
	wire _T_1105 = io_in_d_bits_size == size_1;
	wire _T_1113 = io_in_d_bits_sink == sink;
	wire _T_1117 = io_in_d_bits_denied == denied;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [7:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_72 = {12'd0, inflight_opcodes};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_72 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [15:0] _GEN_74 = {8'd0, inflight_sizes};
	wire [15:0] _a_size_lookup_T_6 = _GEN_74 & _a_size_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_1123 = io_in_a_valid & a_first_1;
	wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source;
	wire [1:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire _T_1126 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [2:0] _GEN_76 = {io_in_a_bits_source, 2'h0};
	wire [3:0] _a_opcodes_set_T = {1'd0, _GEN_76};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _GEN_1 = {15'd0, a_opcodes_set_interm};
	wire [18:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [19:0] _GEN_2 = {15'd0, a_sizes_set_interm};
	wire [19:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire _T_1130 = ~(inflight >> io_in_a_bits_source);
	wire [1:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire [18:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [19:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 20'h00000);
	wire _T_1134 = io_in_d_valid & d_first_1;
	wire _T_1136 = ~_T_930;
	wire _T_1137 = (io_in_d_valid & d_first_1) & ~_T_930;
	wire [1:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_930 ? 2'h1 : 2'h0);
	wire [30:0] _d_opcodes_clr_T_5 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_sizes_clr_T_5 = {15'd0, _a_size_lookup_T_5};
	wire [1:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_1136 ? 2'h1 : 2'h0);
	wire [30:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1136 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [30:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1136 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire same_cycle_resp = _T_1123 & _source_ok_T;
	wire _T_1149 = inflight | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1154 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1155 = (io_in_d_bits_opcode == _GEN_32) | _T_1154;
	wire _T_1159 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1166 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1167 = (io_in_d_bits_opcode == _GEN_48) | _T_1166;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_77 = {4'd0, io_in_d_bits_size};
	wire _T_1171 = _GEN_77 == a_size_lookup;
	wire _T_1181 = (((_T_1134 & a_first_1) & io_in_a_valid) & _source_ok_T) & _T_1136;
	wire _T_1183 = ~io_in_d_ready | io_in_a_ready;
	wire a_set_wo_ready = _GEN_15[0];
	wire d_clr_wo_ready = _GEN_21[0];
	wire _T_1190 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire a_set = _GEN_16[0];
	wire d_clr = _GEN_22[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [7:0] a_sizes_set = _GEN_20[7:0];
	wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [7:0] d_sizes_clr = _GEN_24[7:0];
	wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1199 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [7:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [15:0] _GEN_80 = {8'd0, inflight_sizes_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_80 & _a_size_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_1225 = (io_in_d_valid & d_first_2) & _T_930;
	wire [30:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_930 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1243 = _GEN_77 == c_size_lookup;
	wire [7:0] d_sizes_clr_1 = _GEN_69[7:0];
	wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 8'h00;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 8'h00;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module TLMonitor_1 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_1 = ~io_in_a_bits_source;
	wire source_ok = io_in_a_bits_source | _source_ok_T_1;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_24 = io_in_a_bits_opcode == 3'h6;
	wire _T_26 = io_in_a_bits_size <= 4'hc;
	wire _T_31 = _T_26 & source_ok;
	wire [32:0] _T_37 = $signed(_T_7) & -33'sh000005000;
	wire _T_38 = $signed(_T_37) == 33'sh000000000;
	wire [31:0] _T_39 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_40 = {1'b0, $signed(_T_39)};
	wire [32:0] _T_42 = $signed(_T_40) & -33'sh000001000;
	wire _T_43 = $signed(_T_42) == 33'sh000000000;
	wire [31:0] _T_44 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_45 = {1'b0, $signed(_T_44)};
	wire [32:0] _T_47 = $signed(_T_45) & -33'sh000010000;
	wire _T_48 = $signed(_T_47) == 33'sh000000000;
	wire [31:0] _T_49 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_50 = {1'b0, $signed(_T_49)};
	wire [32:0] _T_52 = $signed(_T_50) & -33'sh000010000;
	wire _T_53 = $signed(_T_52) == 33'sh000000000;
	wire [31:0] _T_54 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_55 = {1'b0, $signed(_T_54)};
	wire [32:0] _T_57 = $signed(_T_55) & -33'sh000011000;
	wire _T_58 = $signed(_T_57) == 33'sh000000000;
	wire [31:0] _T_59 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_60 = {1'b0, $signed(_T_59)};
	wire [32:0] _T_62 = $signed(_T_60) & -33'sh000010000;
	wire _T_63 = $signed(_T_62) == 33'sh000000000;
	wire [31:0] _T_64 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_65 = {1'b0, $signed(_T_64)};
	wire [32:0] _T_67 = $signed(_T_65) & -33'sh004000000;
	wire _T_68 = $signed(_T_67) == 33'sh000000000;
	wire [31:0] _T_69 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_70 = {1'b0, $signed(_T_69)};
	wire [32:0] _T_72 = $signed(_T_70) & -33'sh000001000;
	wire _T_73 = $signed(_T_72) == 33'sh000000000;
	wire [31:0] _T_74 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_75 = {1'b0, $signed(_T_74)};
	wire [32:0] _T_77 = $signed(_T_75) & -33'sh000001000;
	wire _T_78 = $signed(_T_77) == 33'sh000000000;
	wire [31:0] _T_79 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_80 = {1'b0, $signed(_T_79)};
	wire [32:0] _T_82 = $signed(_T_80) & -33'sh000004000;
	wire _T_83 = $signed(_T_82) == 33'sh000000000;
	wire _T_178 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_182 = ~io_in_a_bits_mask;
	wire _T_183 = _T_182 == 4'h0;
	wire _T_187 = ~io_in_a_bits_corrupt;
	wire _T_191 = io_in_a_bits_opcode == 3'h7;
	wire _T_349 = io_in_a_bits_param != 3'h0;
	wire _T_362 = io_in_a_bits_opcode == 3'h4;
	wire _T_383 = _T_26 & _T_43;
	wire _T_385 = io_in_a_bits_size <= 4'h6;
	wire _T_440 = (((((((_T_38 | _T_48) | _T_53) | _T_58) | _T_63) | _T_68) | _T_73) | _T_78) | _T_83;
	wire _T_441 = _T_385 & _T_440;
	wire _T_443 = _T_383 | _T_441;
	wire _T_453 = io_in_a_bits_param == 3'h0;
	wire _T_457 = io_in_a_bits_mask == mask;
	wire _T_465 = io_in_a_bits_opcode == 3'h0;
	wire _T_528 = (((((_T_38 | _T_58) | _T_63) | _T_68) | _T_73) | _T_78) | _T_83;
	wire _T_529 = _T_385 & _T_528;
	wire _T_544 = _T_383 | _T_529;
	wire _T_546 = _T_31 & _T_544;
	wire _T_564 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_659 = ~mask;
	wire [3:0] _T_660 = io_in_a_bits_mask & _T_659;
	wire _T_661 = _T_660 == 4'h0;
	wire _T_665 = io_in_a_bits_opcode == 3'h2;
	wire _T_675 = io_in_a_bits_size <= 4'h2;
	wire _T_724 = ((((((_T_38 | _T_43) | _T_58) | _T_63) | _T_68) | _T_73) | _T_78) | _T_83;
	wire _T_725 = _T_675 & _T_724;
	wire _T_741 = _T_31 & _T_725;
	wire _T_751 = io_in_a_bits_param <= 3'h4;
	wire _T_759 = io_in_a_bits_opcode == 3'h3;
	wire _T_845 = io_in_a_bits_param <= 3'h3;
	wire _T_853 = io_in_a_bits_opcode == 3'h5;
	wire _T_929 = _T_31 & _T_383;
	wire _T_939 = io_in_a_bits_param <= 3'h1;
	wire _T_951 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_3 = ~io_in_d_bits_source;
	wire source_ok_1 = io_in_d_bits_source | _source_ok_T_3;
	wire _T_955 = io_in_d_bits_opcode == 3'h6;
	wire _T_959 = io_in_d_bits_size >= 4'h2;
	wire _T_963 = io_in_d_bits_param == 2'h0;
	wire _T_967 = ~io_in_d_bits_corrupt;
	wire _T_971 = ~io_in_d_bits_denied;
	wire _T_975 = io_in_d_bits_opcode == 3'h4;
	wire _T_986 = io_in_d_bits_param <= 2'h2;
	wire _T_990 = io_in_d_bits_param != 2'h2;
	wire _T_1003 = io_in_d_bits_opcode == 3'h5;
	wire _T_1023 = _T_971 | io_in_d_bits_corrupt;
	wire _T_1032 = io_in_d_bits_opcode == 3'h0;
	wire _T_1049 = io_in_d_bits_opcode == 3'h1;
	wire _T_1067 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg source;
	reg [31:0] address;
	wire _T_1097 = io_in_a_valid & ~a_first;
	wire _T_1098 = io_in_a_bits_opcode == opcode;
	wire _T_1102 = io_in_a_bits_param == param;
	wire _T_1106 = io_in_a_bits_size == size;
	wire _T_1110 = io_in_a_bits_source == source;
	wire _T_1114 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg source_1;
	reg sink;
	reg denied;
	wire _T_1121 = io_in_d_valid & ~d_first;
	wire _T_1122 = io_in_d_bits_opcode == opcode_1;
	wire _T_1126 = io_in_d_bits_param == param_1;
	wire _T_1130 = io_in_d_bits_size == size_1;
	wire _T_1134 = io_in_d_bits_source == source_1;
	wire _T_1138 = io_in_d_bits_sink == sink;
	wire _T_1142 = io_in_d_bits_denied == denied;
	reg [1:0] inflight;
	reg [7:0] inflight_opcodes;
	reg [15:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [3:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [7:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_73 = {8'd0, _a_opcode_lookup_T_1};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0};
	wire [15:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T;
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [15:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _a_size_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_1148 = io_in_a_valid & a_first_1;
	wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source;
	wire [1:0] a_set_wo_ready = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire _T_1151 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [2:0] _GEN_76 = {io_in_a_bits_source, 2'h0};
	wire [3:0] _a_opcodes_set_T = {1'd0, _GEN_76};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _GEN_1 = {15'd0, a_opcodes_set_interm};
	wire [18:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [19:0] _GEN_2 = {15'd0, a_sizes_set_interm};
	wire [19:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire [1:0] _T_1153 = inflight >> io_in_a_bits_source;
	wire _T_1155 = ~_T_1153[0];
	wire [1:0] a_set = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire [18:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [19:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 20'h00000);
	wire _T_1159 = io_in_d_valid & d_first_1;
	wire _T_1161 = ~_T_955;
	wire _T_1162 = (io_in_d_valid & d_first_1) & ~_T_955;
	wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source;
	wire [1:0] d_clr_wo_ready = ((io_in_d_valid & d_first_1) & ~_T_955 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_3 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [30:0] _GEN_4 = {15'd0, _a_size_lookup_T_5};
	wire [30:0] _d_sizes_clr_T_5 = _GEN_4 << _a_size_lookup_T;
	wire [1:0] d_clr = ((_d_first_T & d_first_1) & _T_1161 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1161 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [30:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1161 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_1148 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [1:0] _T_1172 = inflight >> io_in_d_bits_source;
	wire _T_1174 = _T_1172[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1179 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1180 = (io_in_d_bits_opcode == _GEN_32) | _T_1179;
	wire _T_1184 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1191 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1192 = (io_in_d_bits_opcode == _GEN_48) | _T_1191;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_78 = {4'd0, io_in_d_bits_size};
	wire _T_1196 = _GEN_78 == a_size_lookup;
	wire _T_1206 = (((_T_1159 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_1161;
	wire _T_1208 = ~io_in_d_ready | io_in_a_ready;
	wire _T_1215 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [1:0] _inflight_T = inflight | a_set;
	wire [1:0] _inflight_T_1 = ~d_clr;
	wire [1:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [7:0] a_opcodes_set = _GEN_19[7:0];
	wire [7:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [7:0] d_opcodes_clr = _GEN_23[7:0];
	wire [7:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [7:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [15:0] a_sizes_set = _GEN_20[15:0];
	wire [15:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [15:0] d_sizes_clr = _GEN_24[15:0];
	wire [15:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [15:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1224 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [1:0] inflight_1;
	reg [15:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [15:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T;
	wire [15:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _a_size_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_1250 = (io_in_d_valid & d_first_2) & _T_955;
	wire [1:0] d_clr_1 = ((_d_first_T & d_first_2) & _T_955 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_955 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire [1:0] _T_1258 = inflight_1 >> io_in_d_bits_source;
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1268 = _GEN_78 == c_size_lookup;
	wire [1:0] _inflight_T_4 = ~d_clr_1;
	wire [1:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [15:0] d_sizes_clr_1 = _GEN_69[15:0];
	wire [15:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [15:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	reg [31:0] watchdog_1;
	wire _T_1293 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 2'h0;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 8'h00;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 16'h0000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 2'h0;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 16'h0000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLXbar (
	clock,
	reset,
	auto_in_1_a_ready,
	auto_in_1_a_valid,
	auto_in_1_a_bits_opcode,
	auto_in_1_a_bits_param,
	auto_in_1_a_bits_size,
	auto_in_1_a_bits_source,
	auto_in_1_a_bits_address,
	auto_in_1_a_bits_mask,
	auto_in_1_a_bits_data,
	auto_in_1_a_bits_corrupt,
	auto_in_1_d_ready,
	auto_in_1_d_valid,
	auto_in_1_d_bits_opcode,
	auto_in_1_d_bits_param,
	auto_in_1_d_bits_size,
	auto_in_1_d_bits_source,
	auto_in_1_d_bits_sink,
	auto_in_1_d_bits_denied,
	auto_in_1_d_bits_data,
	auto_in_1_d_bits_corrupt,
	auto_in_0_a_ready,
	auto_in_0_a_valid,
	auto_in_0_a_bits_opcode,
	auto_in_0_a_bits_param,
	auto_in_0_a_bits_size,
	auto_in_0_a_bits_source,
	auto_in_0_a_bits_address,
	auto_in_0_a_bits_mask,
	auto_in_0_a_bits_data,
	auto_in_0_a_bits_corrupt,
	auto_in_0_d_ready,
	auto_in_0_d_valid,
	auto_in_0_d_bits_opcode,
	auto_in_0_d_bits_param,
	auto_in_0_d_bits_size,
	auto_in_0_d_bits_sink,
	auto_in_0_d_bits_denied,
	auto_in_0_d_bits_data,
	auto_in_0_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_1_a_ready;
	input auto_in_1_a_valid;
	input [2:0] auto_in_1_a_bits_opcode;
	input [2:0] auto_in_1_a_bits_param;
	input [3:0] auto_in_1_a_bits_size;
	input auto_in_1_a_bits_source;
	input [31:0] auto_in_1_a_bits_address;
	input [3:0] auto_in_1_a_bits_mask;
	input [31:0] auto_in_1_a_bits_data;
	input auto_in_1_a_bits_corrupt;
	input auto_in_1_d_ready;
	output wire auto_in_1_d_valid;
	output wire [2:0] auto_in_1_d_bits_opcode;
	output wire [1:0] auto_in_1_d_bits_param;
	output wire [3:0] auto_in_1_d_bits_size;
	output wire auto_in_1_d_bits_source;
	output wire auto_in_1_d_bits_sink;
	output wire auto_in_1_d_bits_denied;
	output wire [31:0] auto_in_1_d_bits_data;
	output wire auto_in_1_d_bits_corrupt;
	output wire auto_in_0_a_ready;
	input auto_in_0_a_valid;
	input [2:0] auto_in_0_a_bits_opcode;
	input [2:0] auto_in_0_a_bits_param;
	input [3:0] auto_in_0_a_bits_size;
	input auto_in_0_a_bits_source;
	input [31:0] auto_in_0_a_bits_address;
	input [3:0] auto_in_0_a_bits_mask;
	input [31:0] auto_in_0_a_bits_data;
	input auto_in_0_a_bits_corrupt;
	input auto_in_0_d_ready;
	output wire auto_in_0_d_valid;
	output wire [2:0] auto_in_0_d_bits_opcode;
	output wire [1:0] auto_in_0_d_bits_param;
	output wire [3:0] auto_in_0_d_bits_size;
	output wire auto_in_0_d_bits_sink;
	output wire auto_in_0_d_bits_denied;
	output wire [31:0] auto_in_0_d_bits_data;
	output wire auto_in_0_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire [1:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input [1:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire monitor_io_in_a_bits_source;
	wire [31:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [3:0] monitor_io_in_d_bits_size;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire monitor_1_clock;
	wire monitor_1_reset;
	wire monitor_1_io_in_a_ready;
	wire monitor_1_io_in_a_valid;
	wire [2:0] monitor_1_io_in_a_bits_opcode;
	wire [2:0] monitor_1_io_in_a_bits_param;
	wire [3:0] monitor_1_io_in_a_bits_size;
	wire monitor_1_io_in_a_bits_source;
	wire [31:0] monitor_1_io_in_a_bits_address;
	wire [3:0] monitor_1_io_in_a_bits_mask;
	wire monitor_1_io_in_a_bits_corrupt;
	wire monitor_1_io_in_d_ready;
	wire monitor_1_io_in_d_valid;
	wire [2:0] monitor_1_io_in_d_bits_opcode;
	wire [1:0] monitor_1_io_in_d_bits_param;
	wire [3:0] monitor_1_io_in_d_bits_size;
	wire monitor_1_io_in_d_bits_source;
	wire monitor_1_io_in_d_bits_sink;
	wire monitor_1_io_in_d_bits_denied;
	wire monitor_1_io_in_d_bits_corrupt;
	wire [1:0] _GEN_1 = {1'd0, auto_in_0_a_bits_source};
	wire [1:0] in_0_a_bits_source = _GEN_1 | 2'h2;
	wire requestDOI_0_0 = auto_out_d_bits_source == 2'h2;
	wire requestDOI_0_1 = ~auto_out_d_bits_source[1];
	wire [26:0] _beatsAI_decode_T_1 = 27'h0000fff << auto_in_0_a_bits_size;
	wire [11:0] _beatsAI_decode_T_3 = ~_beatsAI_decode_T_1[11:0];
	wire [9:0] beatsAI_decode = _beatsAI_decode_T_3[11:2];
	wire beatsAI_opdata = ~auto_in_0_a_bits_opcode[2];
	wire [9:0] beatsAI_0 = (beatsAI_opdata ? beatsAI_decode : 10'h000);
	wire [26:0] _beatsAI_decode_T_5 = 27'h0000fff << auto_in_1_a_bits_size;
	wire [11:0] _beatsAI_decode_T_7 = ~_beatsAI_decode_T_5[11:0];
	wire [9:0] beatsAI_decode_1 = _beatsAI_decode_T_7[11:2];
	wire beatsAI_opdata_1 = ~auto_in_1_a_bits_opcode[2];
	wire [9:0] beatsAI_1 = (beatsAI_opdata_1 ? beatsAI_decode_1 : 10'h000);
	reg [9:0] beatsLeft;
	wire idle = beatsLeft == 10'h000;
	wire latch = idle & auto_out_a_ready;
	wire [1:0] readys_valid = {auto_in_1_a_valid, auto_in_0_a_valid};
	wire _readys_T_3 = ~reset;
	reg [1:0] readys_mask;
	wire [1:0] _readys_filter_T = ~readys_mask;
	wire [1:0] _readys_filter_T_1 = readys_valid & _readys_filter_T;
	wire [3:0] readys_filter = {_readys_filter_T_1, auto_in_1_a_valid, auto_in_0_a_valid};
	wire [3:0] _GEN_2 = {1'd0, readys_filter[3:1]};
	wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_2;
	wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0};
	wire [3:0] _GEN_3 = {1'd0, _readys_unready_T_1[3:1]};
	wire [3:0] readys_unready = _GEN_3 | _readys_unready_T_4;
	wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0];
	wire [1:0] readys_readys = ~_readys_readys_T_2;
	wire [1:0] _readys_mask_T = readys_readys & readys_valid;
	wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0};
	wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0];
	wire readys_0 = readys_readys[0];
	wire readys_1 = readys_readys[1];
	wire earlyWinner_0 = readys_0 & auto_in_0_a_valid;
	wire earlyWinner_1 = readys_1 & auto_in_1_a_valid;
	wire _prefixOR_T = earlyWinner_0 | earlyWinner_1;
	wire _T_10 = auto_in_0_a_valid | auto_in_1_a_valid;
	wire _T_11 = ~(auto_in_0_a_valid | auto_in_1_a_valid);
	wire [9:0] maskedBeats_0 = (earlyWinner_0 ? beatsAI_0 : 10'h000);
	wire [9:0] maskedBeats_1 = (earlyWinner_1 ? beatsAI_1 : 10'h000);
	wire [9:0] initBeats = maskedBeats_0 | maskedBeats_1;
	reg state_0;
	wire muxStateEarly_0 = (idle ? earlyWinner_0 : state_0);
	reg state_1;
	wire muxStateEarly_1 = (idle ? earlyWinner_1 : state_1);
	wire _out_0_a_earlyValid_T_3 = (state_0 & auto_in_0_a_valid) | (state_1 & auto_in_1_a_valid);
	wire out_2_0_a_earlyValid = (idle ? _T_10 : _out_0_a_earlyValid_T_3);
	wire _beatsLeft_T_2 = auto_out_a_ready & out_2_0_a_earlyValid;
	wire [9:0] _GEN_4 = {9'd0, _beatsLeft_T_2};
	wire [9:0] _beatsLeft_T_4 = beatsLeft - _GEN_4;
	wire allowed_0 = (idle ? readys_0 : state_0);
	wire allowed_1 = (idle ? readys_1 : state_1);
	wire [31:0] _T_27 = (muxStateEarly_0 ? auto_in_0_a_bits_data : 32'h00000000);
	wire [31:0] _T_28 = (muxStateEarly_1 ? auto_in_1_a_bits_data : 32'h00000000);
	wire [3:0] _T_30 = (muxStateEarly_0 ? auto_in_0_a_bits_mask : 4'h0);
	wire [3:0] _T_31 = (muxStateEarly_1 ? auto_in_1_a_bits_mask : 4'h0);
	wire [31:0] _T_33 = (muxStateEarly_0 ? auto_in_0_a_bits_address : 32'h00000000);
	wire [31:0] _T_34 = (muxStateEarly_1 ? auto_in_1_a_bits_address : 32'h00000000);
	wire [1:0] _T_36 = (muxStateEarly_0 ? in_0_a_bits_source : 2'h0);
	wire [1:0] in_1_a_bits_source = {1'd0, auto_in_1_a_bits_source};
	wire [1:0] _T_37 = (muxStateEarly_1 ? in_1_a_bits_source : 2'h0);
	wire [3:0] _T_39 = (muxStateEarly_0 ? auto_in_0_a_bits_size : 4'h0);
	wire [3:0] _T_40 = (muxStateEarly_1 ? auto_in_1_a_bits_size : 4'h0);
	wire [2:0] _T_42 = (muxStateEarly_0 ? auto_in_0_a_bits_param : 3'h0);
	wire [2:0] _T_43 = (muxStateEarly_1 ? auto_in_1_a_bits_param : 3'h0);
	wire [2:0] _T_45 = (muxStateEarly_0 ? auto_in_0_a_bits_opcode : 3'h0);
	wire [2:0] _T_46 = (muxStateEarly_1 ? auto_in_1_a_bits_opcode : 3'h0);
	TLMonitor monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	TLMonitor_1 monitor_1(
		.clock(monitor_1_clock),
		.reset(monitor_1_reset),
		.io_in_a_ready(monitor_1_io_in_a_ready),
		.io_in_a_valid(monitor_1_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_1_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_1_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_1_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_1_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_1_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_1_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_1_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_1_io_in_d_ready),
		.io_in_d_valid(monitor_1_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_1_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_1_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_1_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_1_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_1_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_1_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_1_io_in_d_bits_corrupt)
	);
	assign auto_in_1_a_ready = auto_out_a_ready & allowed_1;
	assign auto_in_1_d_valid = auto_out_d_valid & requestDOI_0_1;
	assign auto_in_1_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_1_d_bits_param = auto_out_d_bits_param;
	assign auto_in_1_d_bits_size = auto_out_d_bits_size;
	assign auto_in_1_d_bits_source = auto_out_d_bits_source[0];
	assign auto_in_1_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_1_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_1_d_bits_data = auto_out_d_bits_data;
	assign auto_in_1_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_in_0_a_ready = auto_out_a_ready & allowed_0;
	assign auto_in_0_d_valid = auto_out_d_valid & requestDOI_0_0;
	assign auto_in_0_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_0_d_bits_param = auto_out_d_bits_param;
	assign auto_in_0_d_bits_size = auto_out_d_bits_size;
	assign auto_in_0_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_0_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_0_d_bits_data = auto_out_d_bits_data;
	assign auto_in_0_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = (idle ? _T_10 : _out_0_a_earlyValid_T_3);
	assign auto_out_a_bits_opcode = _T_45 | _T_46;
	assign auto_out_a_bits_param = _T_42 | _T_43;
	assign auto_out_a_bits_size = _T_39 | _T_40;
	assign auto_out_a_bits_source = _T_36 | _T_37;
	assign auto_out_a_bits_address = _T_33 | _T_34;
	assign auto_out_a_bits_mask = _T_30 | _T_31;
	assign auto_out_a_bits_data = _T_27 | _T_28;
	assign auto_out_a_bits_corrupt = (muxStateEarly_0 & auto_in_0_a_bits_corrupt) | (muxStateEarly_1 & auto_in_1_a_bits_corrupt);
	assign auto_out_d_ready = (requestDOI_0_0 & auto_in_0_d_ready) | (requestDOI_0_1 & auto_in_1_d_ready);
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_out_a_ready & allowed_0;
	assign monitor_io_in_a_valid = auto_in_0_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_0_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_0_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_0_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_0_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_0_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_0_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_0_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_0_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid & requestDOI_0_0;
	assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_io_in_d_bits_param = auto_out_d_bits_param;
	assign monitor_io_in_d_bits_size = auto_out_d_bits_size;
	assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink;
	assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied;
	assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign monitor_1_clock = clock;
	assign monitor_1_reset = reset;
	assign monitor_1_io_in_a_ready = auto_out_a_ready & allowed_1;
	assign monitor_1_io_in_a_valid = auto_in_1_a_valid;
	assign monitor_1_io_in_a_bits_opcode = auto_in_1_a_bits_opcode;
	assign monitor_1_io_in_a_bits_param = auto_in_1_a_bits_param;
	assign monitor_1_io_in_a_bits_size = auto_in_1_a_bits_size;
	assign monitor_1_io_in_a_bits_source = auto_in_1_a_bits_source;
	assign monitor_1_io_in_a_bits_address = auto_in_1_a_bits_address;
	assign monitor_1_io_in_a_bits_mask = auto_in_1_a_bits_mask;
	assign monitor_1_io_in_a_bits_corrupt = auto_in_1_a_bits_corrupt;
	assign monitor_1_io_in_d_ready = auto_in_1_d_ready;
	assign monitor_1_io_in_d_valid = auto_out_d_valid & requestDOI_0_1;
	assign monitor_1_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_1_io_in_d_bits_param = auto_out_d_bits_param;
	assign monitor_1_io_in_d_bits_size = auto_out_d_bits_size;
	assign monitor_1_io_in_d_bits_source = auto_out_d_bits_source[0];
	assign monitor_1_io_in_d_bits_sink = auto_out_d_bits_sink;
	assign monitor_1_io_in_d_bits_denied = auto_out_d_bits_denied;
	assign monitor_1_io_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	always @(posedge clock) begin
		if (reset)
			beatsLeft <= 10'h000;
		else if (latch)
			beatsLeft <= initBeats;
		else
			beatsLeft <= _beatsLeft_T_4;
		if (reset)
			readys_mask <= 2'h3;
		else if (latch & |readys_valid)
			readys_mask <= _readys_mask_T_3;
		if (reset)
			state_0 <= 1'h0;
		else if (idle)
			state_0 <= earlyWinner_0;
		if (reset)
			state_1 <= 1'h0;
		else if (idle)
			state_1 <= earlyWinner_1;
	end
endmodule
module TLMonitor_2 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = ~io_in_a_bits_source;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_5 = ~_source_ok_T;
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_15 = io_in_a_bits_opcode == 3'h6;
	wire _T_17 = io_in_a_bits_size <= 4'hc;
	wire _T_20 = _T_17 & _source_ok_T;
	wire [32:0] _T_26 = $signed(_T_7) & -33'sh000005000;
	wire _T_27 = $signed(_T_26) == 33'sh000000000;
	wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_29 = {1'b0, $signed(_T_28)};
	wire [32:0] _T_31 = $signed(_T_29) & -33'sh000001000;
	wire _T_32 = $signed(_T_31) == 33'sh000000000;
	wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [32:0] _T_36 = $signed(_T_34) & -33'sh000010000;
	wire _T_37 = $signed(_T_36) == 33'sh000000000;
	wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_39 = {1'b0, $signed(_T_38)};
	wire [32:0] _T_41 = $signed(_T_39) & -33'sh000010000;
	wire _T_42 = $signed(_T_41) == 33'sh000000000;
	wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_44 = {1'b0, $signed(_T_43)};
	wire [32:0] _T_46 = $signed(_T_44) & -33'sh000011000;
	wire _T_47 = $signed(_T_46) == 33'sh000000000;
	wire [31:0] _T_48 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_49 = {1'b0, $signed(_T_48)};
	wire [32:0] _T_51 = $signed(_T_49) & -33'sh000010000;
	wire _T_52 = $signed(_T_51) == 33'sh000000000;
	wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_54 = {1'b0, $signed(_T_53)};
	wire [32:0] _T_56 = $signed(_T_54) & -33'sh004000000;
	wire _T_57 = $signed(_T_56) == 33'sh000000000;
	wire [31:0] _T_58 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_59 = {1'b0, $signed(_T_58)};
	wire [32:0] _T_61 = $signed(_T_59) & -33'sh000001000;
	wire _T_62 = $signed(_T_61) == 33'sh000000000;
	wire [31:0] _T_63 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_64 = {1'b0, $signed(_T_63)};
	wire [32:0] _T_66 = $signed(_T_64) & -33'sh000001000;
	wire _T_67 = $signed(_T_66) == 33'sh000000000;
	wire [31:0] _T_68 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_69 = {1'b0, $signed(_T_68)};
	wire [32:0] _T_71 = $signed(_T_69) & -33'sh000004000;
	wire _T_72 = $signed(_T_71) == 33'sh000000000;
	wire _T_167 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_171 = ~io_in_a_bits_mask;
	wire _T_172 = _T_171 == 4'h0;
	wire _T_176 = ~io_in_a_bits_corrupt;
	wire _T_180 = io_in_a_bits_opcode == 3'h7;
	wire _T_336 = io_in_a_bits_param != 3'h0;
	wire _T_349 = io_in_a_bits_opcode == 3'h4;
	wire _T_368 = _T_17 & _T_32;
	wire _T_370 = io_in_a_bits_size <= 4'h6;
	wire _T_425 = (((((((_T_27 | _T_37) | _T_42) | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_426 = _T_370 & _T_425;
	wire _T_428 = _T_368 | _T_426;
	wire _T_438 = io_in_a_bits_param == 3'h0;
	wire _T_442 = io_in_a_bits_mask == mask;
	wire _T_450 = io_in_a_bits_opcode == 3'h0;
	wire _T_511 = (((((_T_27 | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_512 = _T_370 & _T_511;
	wire _T_527 = _T_368 | _T_512;
	wire _T_529 = _T_20 & _T_527;
	wire _T_547 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_640 = ~mask;
	wire [3:0] _T_641 = io_in_a_bits_mask & _T_640;
	wire _T_642 = _T_641 == 4'h0;
	wire _T_646 = io_in_a_bits_opcode == 3'h2;
	wire _T_654 = io_in_a_bits_size <= 4'h2;
	wire _T_703 = ((((((_T_27 | _T_32) | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_704 = _T_654 & _T_703;
	wire _T_720 = _T_20 & _T_704;
	wire _T_730 = io_in_a_bits_param <= 3'h4;
	wire _T_738 = io_in_a_bits_opcode == 3'h3;
	wire _T_822 = io_in_a_bits_param <= 3'h3;
	wire _T_830 = io_in_a_bits_opcode == 3'h5;
	wire _T_904 = _T_20 & _T_368;
	wire _T_914 = io_in_a_bits_param <= 3'h1;
	wire _T_926 = io_in_d_bits_opcode <= 3'h6;
	wire _T_930 = io_in_d_bits_opcode == 3'h6;
	wire _T_934 = io_in_d_bits_size >= 4'h2;
	wire _T_938 = io_in_d_bits_param == 2'h0;
	wire _T_942 = ~io_in_d_bits_corrupt;
	wire _T_946 = ~io_in_d_bits_denied;
	wire _T_950 = io_in_d_bits_opcode == 3'h4;
	wire _T_961 = io_in_d_bits_param <= 2'h2;
	wire _T_965 = io_in_d_bits_param != 2'h2;
	wire _T_978 = io_in_d_bits_opcode == 3'h5;
	wire _T_998 = _T_946 | io_in_d_bits_corrupt;
	wire _T_1007 = io_in_d_bits_opcode == 3'h0;
	wire _T_1024 = io_in_d_bits_opcode == 3'h1;
	wire _T_1042 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg source;
	reg [31:0] address;
	wire _T_1072 = io_in_a_valid & ~a_first;
	wire _T_1073 = io_in_a_bits_opcode == opcode;
	wire _T_1077 = io_in_a_bits_param == param;
	wire _T_1081 = io_in_a_bits_size == size;
	wire _T_1085 = io_in_a_bits_source == source;
	wire _T_1089 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg sink;
	reg denied;
	wire _T_1096 = io_in_d_valid & ~d_first;
	wire _T_1097 = io_in_d_bits_opcode == opcode_1;
	wire _T_1101 = io_in_d_bits_param == param_1;
	wire _T_1105 = io_in_d_bits_size == size_1;
	wire _T_1113 = io_in_d_bits_sink == sink;
	wire _T_1117 = io_in_d_bits_denied == denied;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [7:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_72 = {12'd0, inflight_opcodes};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_72 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [15:0] _GEN_74 = {8'd0, inflight_sizes};
	wire [15:0] _a_size_lookup_T_6 = _GEN_74 & _a_size_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_1123 = io_in_a_valid & a_first_1;
	wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source;
	wire [1:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire _T_1126 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [2:0] _GEN_76 = {io_in_a_bits_source, 2'h0};
	wire [3:0] _a_opcodes_set_T = {1'd0, _GEN_76};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _GEN_1 = {15'd0, a_opcodes_set_interm};
	wire [18:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [19:0] _GEN_2 = {15'd0, a_sizes_set_interm};
	wire [19:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire _T_1130 = ~(inflight >> io_in_a_bits_source);
	wire [1:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire [18:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [19:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 20'h00000);
	wire _T_1134 = io_in_d_valid & d_first_1;
	wire _T_1136 = ~_T_930;
	wire _T_1137 = (io_in_d_valid & d_first_1) & ~_T_930;
	wire [1:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_930 ? 2'h1 : 2'h0);
	wire [30:0] _d_opcodes_clr_T_5 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_sizes_clr_T_5 = {15'd0, _a_size_lookup_T_5};
	wire [1:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_1136 ? 2'h1 : 2'h0);
	wire [30:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1136 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [30:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1136 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire same_cycle_resp = _T_1123 & _source_ok_T;
	wire _T_1149 = inflight | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1154 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1155 = (io_in_d_bits_opcode == _GEN_32) | _T_1154;
	wire _T_1159 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1166 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1167 = (io_in_d_bits_opcode == _GEN_48) | _T_1166;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_77 = {4'd0, io_in_d_bits_size};
	wire _T_1171 = _GEN_77 == a_size_lookup;
	wire _T_1181 = (((_T_1134 & a_first_1) & io_in_a_valid) & _source_ok_T) & _T_1136;
	wire _T_1183 = ~io_in_d_ready | io_in_a_ready;
	wire a_set_wo_ready = _GEN_15[0];
	wire d_clr_wo_ready = _GEN_21[0];
	wire _T_1190 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire a_set = _GEN_16[0];
	wire d_clr = _GEN_22[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [7:0] a_sizes_set = _GEN_20[7:0];
	wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [7:0] d_sizes_clr = _GEN_24[7:0];
	wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1199 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [7:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [15:0] _GEN_80 = {8'd0, inflight_sizes_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_80 & _a_size_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_1225 = (io_in_d_valid & d_first_2) & _T_930;
	wire [30:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_930 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1243 = _GEN_77 == c_size_lookup;
	wire [7:0] d_sizes_clr_1 = _GEN_69[7:0];
	wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 8'h00;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 8'h00;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module TLMonitor_3 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_1 = ~io_in_a_bits_source;
	wire source_ok = io_in_a_bits_source | _source_ok_T_1;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_24 = io_in_a_bits_opcode == 3'h6;
	wire _T_26 = io_in_a_bits_size <= 4'hc;
	wire _T_31 = _T_26 & source_ok;
	wire [32:0] _T_37 = $signed(_T_7) & -33'sh000005000;
	wire _T_38 = $signed(_T_37) == 33'sh000000000;
	wire [31:0] _T_39 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_40 = {1'b0, $signed(_T_39)};
	wire [32:0] _T_42 = $signed(_T_40) & -33'sh000001000;
	wire _T_43 = $signed(_T_42) == 33'sh000000000;
	wire [31:0] _T_44 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_45 = {1'b0, $signed(_T_44)};
	wire [32:0] _T_47 = $signed(_T_45) & -33'sh000010000;
	wire _T_48 = $signed(_T_47) == 33'sh000000000;
	wire [31:0] _T_49 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_50 = {1'b0, $signed(_T_49)};
	wire [32:0] _T_52 = $signed(_T_50) & -33'sh000010000;
	wire _T_53 = $signed(_T_52) == 33'sh000000000;
	wire [31:0] _T_54 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_55 = {1'b0, $signed(_T_54)};
	wire [32:0] _T_57 = $signed(_T_55) & -33'sh000011000;
	wire _T_58 = $signed(_T_57) == 33'sh000000000;
	wire [31:0] _T_59 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_60 = {1'b0, $signed(_T_59)};
	wire [32:0] _T_62 = $signed(_T_60) & -33'sh000010000;
	wire _T_63 = $signed(_T_62) == 33'sh000000000;
	wire [31:0] _T_64 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_65 = {1'b0, $signed(_T_64)};
	wire [32:0] _T_67 = $signed(_T_65) & -33'sh004000000;
	wire _T_68 = $signed(_T_67) == 33'sh000000000;
	wire [31:0] _T_69 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_70 = {1'b0, $signed(_T_69)};
	wire [32:0] _T_72 = $signed(_T_70) & -33'sh000001000;
	wire _T_73 = $signed(_T_72) == 33'sh000000000;
	wire [31:0] _T_74 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_75 = {1'b0, $signed(_T_74)};
	wire [32:0] _T_77 = $signed(_T_75) & -33'sh000001000;
	wire _T_78 = $signed(_T_77) == 33'sh000000000;
	wire [31:0] _T_79 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_80 = {1'b0, $signed(_T_79)};
	wire [32:0] _T_82 = $signed(_T_80) & -33'sh000004000;
	wire _T_83 = $signed(_T_82) == 33'sh000000000;
	wire _T_178 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_182 = ~io_in_a_bits_mask;
	wire _T_183 = _T_182 == 4'h0;
	wire _T_187 = ~io_in_a_bits_corrupt;
	wire _T_191 = io_in_a_bits_opcode == 3'h7;
	wire _T_349 = io_in_a_bits_param != 3'h0;
	wire _T_362 = io_in_a_bits_opcode == 3'h4;
	wire _T_383 = _T_26 & _T_43;
	wire _T_385 = io_in_a_bits_size <= 4'h6;
	wire _T_440 = (((((((_T_38 | _T_48) | _T_53) | _T_58) | _T_63) | _T_68) | _T_73) | _T_78) | _T_83;
	wire _T_441 = _T_385 & _T_440;
	wire _T_443 = _T_383 | _T_441;
	wire _T_453 = io_in_a_bits_param == 3'h0;
	wire _T_457 = io_in_a_bits_mask == mask;
	wire _T_465 = io_in_a_bits_opcode == 3'h0;
	wire _T_528 = (((((_T_38 | _T_58) | _T_63) | _T_68) | _T_73) | _T_78) | _T_83;
	wire _T_529 = _T_385 & _T_528;
	wire _T_544 = _T_383 | _T_529;
	wire _T_546 = _T_31 & _T_544;
	wire _T_564 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_659 = ~mask;
	wire [3:0] _T_660 = io_in_a_bits_mask & _T_659;
	wire _T_661 = _T_660 == 4'h0;
	wire _T_665 = io_in_a_bits_opcode == 3'h2;
	wire _T_675 = io_in_a_bits_size <= 4'h2;
	wire _T_724 = ((((((_T_38 | _T_43) | _T_58) | _T_63) | _T_68) | _T_73) | _T_78) | _T_83;
	wire _T_725 = _T_675 & _T_724;
	wire _T_741 = _T_31 & _T_725;
	wire _T_751 = io_in_a_bits_param <= 3'h4;
	wire _T_759 = io_in_a_bits_opcode == 3'h3;
	wire _T_845 = io_in_a_bits_param <= 3'h3;
	wire _T_853 = io_in_a_bits_opcode == 3'h5;
	wire _T_929 = _T_31 & _T_383;
	wire _T_939 = io_in_a_bits_param <= 3'h1;
	wire _T_951 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_3 = ~io_in_d_bits_source;
	wire source_ok_1 = io_in_d_bits_source | _source_ok_T_3;
	wire _T_955 = io_in_d_bits_opcode == 3'h6;
	wire _T_959 = io_in_d_bits_size >= 4'h2;
	wire _T_963 = io_in_d_bits_param == 2'h0;
	wire _T_967 = ~io_in_d_bits_corrupt;
	wire _T_971 = ~io_in_d_bits_denied;
	wire _T_975 = io_in_d_bits_opcode == 3'h4;
	wire _T_986 = io_in_d_bits_param <= 2'h2;
	wire _T_990 = io_in_d_bits_param != 2'h2;
	wire _T_1003 = io_in_d_bits_opcode == 3'h5;
	wire _T_1023 = _T_971 | io_in_d_bits_corrupt;
	wire _T_1032 = io_in_d_bits_opcode == 3'h0;
	wire _T_1049 = io_in_d_bits_opcode == 3'h1;
	wire _T_1067 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg source;
	reg [31:0] address;
	wire _T_1097 = io_in_a_valid & ~a_first;
	wire _T_1098 = io_in_a_bits_opcode == opcode;
	wire _T_1102 = io_in_a_bits_param == param;
	wire _T_1106 = io_in_a_bits_size == size;
	wire _T_1110 = io_in_a_bits_source == source;
	wire _T_1114 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg source_1;
	reg sink;
	reg denied;
	wire _T_1121 = io_in_d_valid & ~d_first;
	wire _T_1122 = io_in_d_bits_opcode == opcode_1;
	wire _T_1126 = io_in_d_bits_param == param_1;
	wire _T_1130 = io_in_d_bits_size == size_1;
	wire _T_1134 = io_in_d_bits_source == source_1;
	wire _T_1138 = io_in_d_bits_sink == sink;
	wire _T_1142 = io_in_d_bits_denied == denied;
	reg [1:0] inflight;
	reg [7:0] inflight_opcodes;
	reg [15:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [3:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [7:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_73 = {8'd0, _a_opcode_lookup_T_1};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0};
	wire [15:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T;
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [15:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _a_size_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_1148 = io_in_a_valid & a_first_1;
	wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source;
	wire [1:0] a_set_wo_ready = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire _T_1151 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [2:0] _GEN_76 = {io_in_a_bits_source, 2'h0};
	wire [3:0] _a_opcodes_set_T = {1'd0, _GEN_76};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _GEN_1 = {15'd0, a_opcodes_set_interm};
	wire [18:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [19:0] _GEN_2 = {15'd0, a_sizes_set_interm};
	wire [19:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire [1:0] _T_1153 = inflight >> io_in_a_bits_source;
	wire _T_1155 = ~_T_1153[0];
	wire [1:0] a_set = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire [18:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [19:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 20'h00000);
	wire _T_1159 = io_in_d_valid & d_first_1;
	wire _T_1161 = ~_T_955;
	wire _T_1162 = (io_in_d_valid & d_first_1) & ~_T_955;
	wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source;
	wire [1:0] d_clr_wo_ready = ((io_in_d_valid & d_first_1) & ~_T_955 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_3 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [30:0] _GEN_4 = {15'd0, _a_size_lookup_T_5};
	wire [30:0] _d_sizes_clr_T_5 = _GEN_4 << _a_size_lookup_T;
	wire [1:0] d_clr = ((_d_first_T & d_first_1) & _T_1161 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1161 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [30:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1161 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_1148 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [1:0] _T_1172 = inflight >> io_in_d_bits_source;
	wire _T_1174 = _T_1172[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1179 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1180 = (io_in_d_bits_opcode == _GEN_32) | _T_1179;
	wire _T_1184 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1191 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1192 = (io_in_d_bits_opcode == _GEN_48) | _T_1191;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_78 = {4'd0, io_in_d_bits_size};
	wire _T_1196 = _GEN_78 == a_size_lookup;
	wire _T_1206 = (((_T_1159 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_1161;
	wire _T_1208 = ~io_in_d_ready | io_in_a_ready;
	wire _T_1215 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [1:0] _inflight_T = inflight | a_set;
	wire [1:0] _inflight_T_1 = ~d_clr;
	wire [1:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [7:0] a_opcodes_set = _GEN_19[7:0];
	wire [7:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [7:0] d_opcodes_clr = _GEN_23[7:0];
	wire [7:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [7:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [15:0] a_sizes_set = _GEN_20[15:0];
	wire [15:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [15:0] d_sizes_clr = _GEN_24[15:0];
	wire [15:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [15:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1224 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [1:0] inflight_1;
	reg [15:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [15:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T;
	wire [15:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _a_size_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_1250 = (io_in_d_valid & d_first_2) & _T_955;
	wire [1:0] d_clr_1 = ((_d_first_T & d_first_2) & _T_955 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_955 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire [1:0] _T_1258 = inflight_1 >> io_in_d_bits_source;
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1268 = _GEN_78 == c_size_lookup;
	wire [1:0] _inflight_T_4 = ~d_clr_1;
	wire [1:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [15:0] d_sizes_clr_1 = _GEN_69[15:0];
	wire [15:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [15:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	reg [31:0] watchdog_1;
	wire _T_1293 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 2'h0;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 8'h00;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 16'h0000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 2'h0;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 16'h0000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLFIFOFixer (
	clock,
	reset,
	auto_in_1_a_ready,
	auto_in_1_a_valid,
	auto_in_1_a_bits_opcode,
	auto_in_1_a_bits_param,
	auto_in_1_a_bits_size,
	auto_in_1_a_bits_source,
	auto_in_1_a_bits_address,
	auto_in_1_a_bits_mask,
	auto_in_1_a_bits_data,
	auto_in_1_a_bits_corrupt,
	auto_in_1_d_ready,
	auto_in_1_d_valid,
	auto_in_1_d_bits_opcode,
	auto_in_1_d_bits_param,
	auto_in_1_d_bits_size,
	auto_in_1_d_bits_source,
	auto_in_1_d_bits_sink,
	auto_in_1_d_bits_denied,
	auto_in_1_d_bits_data,
	auto_in_1_d_bits_corrupt,
	auto_in_0_a_ready,
	auto_in_0_a_valid,
	auto_in_0_a_bits_opcode,
	auto_in_0_a_bits_param,
	auto_in_0_a_bits_size,
	auto_in_0_a_bits_source,
	auto_in_0_a_bits_address,
	auto_in_0_a_bits_mask,
	auto_in_0_a_bits_data,
	auto_in_0_a_bits_corrupt,
	auto_in_0_d_ready,
	auto_in_0_d_valid,
	auto_in_0_d_bits_opcode,
	auto_in_0_d_bits_param,
	auto_in_0_d_bits_size,
	auto_in_0_d_bits_sink,
	auto_in_0_d_bits_denied,
	auto_in_0_d_bits_data,
	auto_in_0_d_bits_corrupt,
	auto_out_1_a_ready,
	auto_out_1_a_valid,
	auto_out_1_a_bits_opcode,
	auto_out_1_a_bits_param,
	auto_out_1_a_bits_size,
	auto_out_1_a_bits_source,
	auto_out_1_a_bits_address,
	auto_out_1_a_bits_mask,
	auto_out_1_a_bits_data,
	auto_out_1_a_bits_corrupt,
	auto_out_1_d_ready,
	auto_out_1_d_valid,
	auto_out_1_d_bits_opcode,
	auto_out_1_d_bits_param,
	auto_out_1_d_bits_size,
	auto_out_1_d_bits_source,
	auto_out_1_d_bits_sink,
	auto_out_1_d_bits_denied,
	auto_out_1_d_bits_data,
	auto_out_1_d_bits_corrupt,
	auto_out_0_a_ready,
	auto_out_0_a_valid,
	auto_out_0_a_bits_opcode,
	auto_out_0_a_bits_param,
	auto_out_0_a_bits_size,
	auto_out_0_a_bits_source,
	auto_out_0_a_bits_address,
	auto_out_0_a_bits_mask,
	auto_out_0_a_bits_data,
	auto_out_0_a_bits_corrupt,
	auto_out_0_d_ready,
	auto_out_0_d_valid,
	auto_out_0_d_bits_opcode,
	auto_out_0_d_bits_param,
	auto_out_0_d_bits_size,
	auto_out_0_d_bits_sink,
	auto_out_0_d_bits_denied,
	auto_out_0_d_bits_data,
	auto_out_0_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_1_a_ready;
	input auto_in_1_a_valid;
	input [2:0] auto_in_1_a_bits_opcode;
	input [2:0] auto_in_1_a_bits_param;
	input [3:0] auto_in_1_a_bits_size;
	input auto_in_1_a_bits_source;
	input [31:0] auto_in_1_a_bits_address;
	input [3:0] auto_in_1_a_bits_mask;
	input [31:0] auto_in_1_a_bits_data;
	input auto_in_1_a_bits_corrupt;
	input auto_in_1_d_ready;
	output wire auto_in_1_d_valid;
	output wire [2:0] auto_in_1_d_bits_opcode;
	output wire [1:0] auto_in_1_d_bits_param;
	output wire [3:0] auto_in_1_d_bits_size;
	output wire auto_in_1_d_bits_source;
	output wire auto_in_1_d_bits_sink;
	output wire auto_in_1_d_bits_denied;
	output wire [31:0] auto_in_1_d_bits_data;
	output wire auto_in_1_d_bits_corrupt;
	output wire auto_in_0_a_ready;
	input auto_in_0_a_valid;
	input [2:0] auto_in_0_a_bits_opcode;
	input [2:0] auto_in_0_a_bits_param;
	input [3:0] auto_in_0_a_bits_size;
	input auto_in_0_a_bits_source;
	input [31:0] auto_in_0_a_bits_address;
	input [3:0] auto_in_0_a_bits_mask;
	input [31:0] auto_in_0_a_bits_data;
	input auto_in_0_a_bits_corrupt;
	input auto_in_0_d_ready;
	output wire auto_in_0_d_valid;
	output wire [2:0] auto_in_0_d_bits_opcode;
	output wire [1:0] auto_in_0_d_bits_param;
	output wire [3:0] auto_in_0_d_bits_size;
	output wire auto_in_0_d_bits_sink;
	output wire auto_in_0_d_bits_denied;
	output wire [31:0] auto_in_0_d_bits_data;
	output wire auto_in_0_d_bits_corrupt;
	input auto_out_1_a_ready;
	output wire auto_out_1_a_valid;
	output wire [2:0] auto_out_1_a_bits_opcode;
	output wire [2:0] auto_out_1_a_bits_param;
	output wire [3:0] auto_out_1_a_bits_size;
	output wire auto_out_1_a_bits_source;
	output wire [31:0] auto_out_1_a_bits_address;
	output wire [3:0] auto_out_1_a_bits_mask;
	output wire [31:0] auto_out_1_a_bits_data;
	output wire auto_out_1_a_bits_corrupt;
	output wire auto_out_1_d_ready;
	input auto_out_1_d_valid;
	input [2:0] auto_out_1_d_bits_opcode;
	input [1:0] auto_out_1_d_bits_param;
	input [3:0] auto_out_1_d_bits_size;
	input auto_out_1_d_bits_source;
	input auto_out_1_d_bits_sink;
	input auto_out_1_d_bits_denied;
	input [31:0] auto_out_1_d_bits_data;
	input auto_out_1_d_bits_corrupt;
	input auto_out_0_a_ready;
	output wire auto_out_0_a_valid;
	output wire [2:0] auto_out_0_a_bits_opcode;
	output wire [2:0] auto_out_0_a_bits_param;
	output wire [3:0] auto_out_0_a_bits_size;
	output wire auto_out_0_a_bits_source;
	output wire [31:0] auto_out_0_a_bits_address;
	output wire [3:0] auto_out_0_a_bits_mask;
	output wire [31:0] auto_out_0_a_bits_data;
	output wire auto_out_0_a_bits_corrupt;
	output wire auto_out_0_d_ready;
	input auto_out_0_d_valid;
	input [2:0] auto_out_0_d_bits_opcode;
	input [1:0] auto_out_0_d_bits_param;
	input [3:0] auto_out_0_d_bits_size;
	input auto_out_0_d_bits_sink;
	input auto_out_0_d_bits_denied;
	input [31:0] auto_out_0_d_bits_data;
	input auto_out_0_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire monitor_io_in_a_bits_source;
	wire [31:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [3:0] monitor_io_in_d_bits_size;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire monitor_1_clock;
	wire monitor_1_reset;
	wire monitor_1_io_in_a_ready;
	wire monitor_1_io_in_a_valid;
	wire [2:0] monitor_1_io_in_a_bits_opcode;
	wire [2:0] monitor_1_io_in_a_bits_param;
	wire [3:0] monitor_1_io_in_a_bits_size;
	wire monitor_1_io_in_a_bits_source;
	wire [31:0] monitor_1_io_in_a_bits_address;
	wire [3:0] monitor_1_io_in_a_bits_mask;
	wire monitor_1_io_in_a_bits_corrupt;
	wire monitor_1_io_in_d_ready;
	wire monitor_1_io_in_d_valid;
	wire [2:0] monitor_1_io_in_d_bits_opcode;
	wire [1:0] monitor_1_io_in_d_bits_param;
	wire [3:0] monitor_1_io_in_d_bits_size;
	wire monitor_1_io_in_d_bits_source;
	wire monitor_1_io_in_d_bits_sink;
	wire monitor_1_io_in_d_bits_denied;
	wire monitor_1_io_in_d_bits_corrupt;
	TLMonitor_2 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	TLMonitor_3 monitor_1(
		.clock(monitor_1_clock),
		.reset(monitor_1_reset),
		.io_in_a_ready(monitor_1_io_in_a_ready),
		.io_in_a_valid(monitor_1_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_1_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_1_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_1_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_1_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_1_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_1_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_1_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_1_io_in_d_ready),
		.io_in_d_valid(monitor_1_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_1_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_1_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_1_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_1_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_1_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_1_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_1_io_in_d_bits_corrupt)
	);
	assign auto_in_1_a_ready = auto_out_1_a_ready;
	assign auto_in_1_d_valid = auto_out_1_d_valid;
	assign auto_in_1_d_bits_opcode = auto_out_1_d_bits_opcode;
	assign auto_in_1_d_bits_param = auto_out_1_d_bits_param;
	assign auto_in_1_d_bits_size = auto_out_1_d_bits_size;
	assign auto_in_1_d_bits_source = auto_out_1_d_bits_source;
	assign auto_in_1_d_bits_sink = auto_out_1_d_bits_sink;
	assign auto_in_1_d_bits_denied = auto_out_1_d_bits_denied;
	assign auto_in_1_d_bits_data = auto_out_1_d_bits_data;
	assign auto_in_1_d_bits_corrupt = auto_out_1_d_bits_corrupt;
	assign auto_in_0_a_ready = auto_out_0_a_ready;
	assign auto_in_0_d_valid = auto_out_0_d_valid;
	assign auto_in_0_d_bits_opcode = auto_out_0_d_bits_opcode;
	assign auto_in_0_d_bits_param = auto_out_0_d_bits_param;
	assign auto_in_0_d_bits_size = auto_out_0_d_bits_size;
	assign auto_in_0_d_bits_sink = auto_out_0_d_bits_sink;
	assign auto_in_0_d_bits_denied = auto_out_0_d_bits_denied;
	assign auto_in_0_d_bits_data = auto_out_0_d_bits_data;
	assign auto_in_0_d_bits_corrupt = auto_out_0_d_bits_corrupt;
	assign auto_out_1_a_valid = auto_in_1_a_valid;
	assign auto_out_1_a_bits_opcode = auto_in_1_a_bits_opcode;
	assign auto_out_1_a_bits_param = auto_in_1_a_bits_param;
	assign auto_out_1_a_bits_size = auto_in_1_a_bits_size;
	assign auto_out_1_a_bits_source = auto_in_1_a_bits_source;
	assign auto_out_1_a_bits_address = auto_in_1_a_bits_address;
	assign auto_out_1_a_bits_mask = auto_in_1_a_bits_mask;
	assign auto_out_1_a_bits_data = auto_in_1_a_bits_data;
	assign auto_out_1_a_bits_corrupt = auto_in_1_a_bits_corrupt;
	assign auto_out_1_d_ready = auto_in_1_d_ready;
	assign auto_out_0_a_valid = auto_in_0_a_valid;
	assign auto_out_0_a_bits_opcode = auto_in_0_a_bits_opcode;
	assign auto_out_0_a_bits_param = auto_in_0_a_bits_param;
	assign auto_out_0_a_bits_size = auto_in_0_a_bits_size;
	assign auto_out_0_a_bits_source = auto_in_0_a_bits_source;
	assign auto_out_0_a_bits_address = auto_in_0_a_bits_address;
	assign auto_out_0_a_bits_mask = auto_in_0_a_bits_mask;
	assign auto_out_0_a_bits_data = auto_in_0_a_bits_data;
	assign auto_out_0_a_bits_corrupt = auto_in_0_a_bits_corrupt;
	assign auto_out_0_d_ready = auto_in_0_d_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_out_0_a_ready;
	assign monitor_io_in_a_valid = auto_in_0_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_0_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_0_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_0_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_0_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_0_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_0_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_0_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_0_d_ready;
	assign monitor_io_in_d_valid = auto_out_0_d_valid;
	assign monitor_io_in_d_bits_opcode = auto_out_0_d_bits_opcode;
	assign monitor_io_in_d_bits_param = auto_out_0_d_bits_param;
	assign monitor_io_in_d_bits_size = auto_out_0_d_bits_size;
	assign monitor_io_in_d_bits_sink = auto_out_0_d_bits_sink;
	assign monitor_io_in_d_bits_denied = auto_out_0_d_bits_denied;
	assign monitor_io_in_d_bits_corrupt = auto_out_0_d_bits_corrupt;
	assign monitor_1_clock = clock;
	assign monitor_1_reset = reset;
	assign monitor_1_io_in_a_ready = auto_out_1_a_ready;
	assign monitor_1_io_in_a_valid = auto_in_1_a_valid;
	assign monitor_1_io_in_a_bits_opcode = auto_in_1_a_bits_opcode;
	assign monitor_1_io_in_a_bits_param = auto_in_1_a_bits_param;
	assign monitor_1_io_in_a_bits_size = auto_in_1_a_bits_size;
	assign monitor_1_io_in_a_bits_source = auto_in_1_a_bits_source;
	assign monitor_1_io_in_a_bits_address = auto_in_1_a_bits_address;
	assign monitor_1_io_in_a_bits_mask = auto_in_1_a_bits_mask;
	assign monitor_1_io_in_a_bits_corrupt = auto_in_1_a_bits_corrupt;
	assign monitor_1_io_in_d_ready = auto_in_1_d_ready;
	assign monitor_1_io_in_d_valid = auto_out_1_d_valid;
	assign monitor_1_io_in_d_bits_opcode = auto_out_1_d_bits_opcode;
	assign monitor_1_io_in_d_bits_param = auto_out_1_d_bits_param;
	assign monitor_1_io_in_d_bits_size = auto_out_1_d_bits_size;
	assign monitor_1_io_in_d_bits_source = auto_out_1_d_bits_source;
	assign monitor_1_io_in_d_bits_sink = auto_out_1_d_bits_sink;
	assign monitor_1_io_in_d_bits_denied = auto_out_1_d_bits_denied;
	assign monitor_1_io_in_d_bits_corrupt = auto_out_1_d_bits_corrupt;
endmodule
module TLWidthWidget (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input [1:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire [1:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire [1:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input [1:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module TLInterconnectCoupler (
	auto_widget_in_a_ready,
	auto_widget_in_a_valid,
	auto_widget_in_a_bits_opcode,
	auto_widget_in_a_bits_param,
	auto_widget_in_a_bits_size,
	auto_widget_in_a_bits_source,
	auto_widget_in_a_bits_address,
	auto_widget_in_a_bits_mask,
	auto_widget_in_a_bits_data,
	auto_widget_in_a_bits_corrupt,
	auto_widget_in_d_ready,
	auto_widget_in_d_valid,
	auto_widget_in_d_bits_opcode,
	auto_widget_in_d_bits_param,
	auto_widget_in_d_bits_size,
	auto_widget_in_d_bits_source,
	auto_widget_in_d_bits_sink,
	auto_widget_in_d_bits_denied,
	auto_widget_in_d_bits_data,
	auto_widget_in_d_bits_corrupt,
	auto_bus_xing_out_a_ready,
	auto_bus_xing_out_a_valid,
	auto_bus_xing_out_a_bits_opcode,
	auto_bus_xing_out_a_bits_param,
	auto_bus_xing_out_a_bits_size,
	auto_bus_xing_out_a_bits_source,
	auto_bus_xing_out_a_bits_address,
	auto_bus_xing_out_a_bits_mask,
	auto_bus_xing_out_a_bits_data,
	auto_bus_xing_out_a_bits_corrupt,
	auto_bus_xing_out_d_ready,
	auto_bus_xing_out_d_valid,
	auto_bus_xing_out_d_bits_opcode,
	auto_bus_xing_out_d_bits_param,
	auto_bus_xing_out_d_bits_size,
	auto_bus_xing_out_d_bits_source,
	auto_bus_xing_out_d_bits_sink,
	auto_bus_xing_out_d_bits_denied,
	auto_bus_xing_out_d_bits_data,
	auto_bus_xing_out_d_bits_corrupt
);
	output wire auto_widget_in_a_ready;
	input auto_widget_in_a_valid;
	input [2:0] auto_widget_in_a_bits_opcode;
	input [2:0] auto_widget_in_a_bits_param;
	input [3:0] auto_widget_in_a_bits_size;
	input [1:0] auto_widget_in_a_bits_source;
	input [31:0] auto_widget_in_a_bits_address;
	input [3:0] auto_widget_in_a_bits_mask;
	input [31:0] auto_widget_in_a_bits_data;
	input auto_widget_in_a_bits_corrupt;
	input auto_widget_in_d_ready;
	output wire auto_widget_in_d_valid;
	output wire [2:0] auto_widget_in_d_bits_opcode;
	output wire [1:0] auto_widget_in_d_bits_param;
	output wire [3:0] auto_widget_in_d_bits_size;
	output wire [1:0] auto_widget_in_d_bits_source;
	output wire auto_widget_in_d_bits_sink;
	output wire auto_widget_in_d_bits_denied;
	output wire [31:0] auto_widget_in_d_bits_data;
	output wire auto_widget_in_d_bits_corrupt;
	input auto_bus_xing_out_a_ready;
	output wire auto_bus_xing_out_a_valid;
	output wire [2:0] auto_bus_xing_out_a_bits_opcode;
	output wire [2:0] auto_bus_xing_out_a_bits_param;
	output wire [3:0] auto_bus_xing_out_a_bits_size;
	output wire [1:0] auto_bus_xing_out_a_bits_source;
	output wire [31:0] auto_bus_xing_out_a_bits_address;
	output wire [3:0] auto_bus_xing_out_a_bits_mask;
	output wire [31:0] auto_bus_xing_out_a_bits_data;
	output wire auto_bus_xing_out_a_bits_corrupt;
	output wire auto_bus_xing_out_d_ready;
	input auto_bus_xing_out_d_valid;
	input [2:0] auto_bus_xing_out_d_bits_opcode;
	input [1:0] auto_bus_xing_out_d_bits_param;
	input [3:0] auto_bus_xing_out_d_bits_size;
	input [1:0] auto_bus_xing_out_d_bits_source;
	input auto_bus_xing_out_d_bits_sink;
	input auto_bus_xing_out_d_bits_denied;
	input [31:0] auto_bus_xing_out_d_bits_data;
	input auto_bus_xing_out_d_bits_corrupt;
	wire widget_auto_in_a_ready;
	wire widget_auto_in_a_valid;
	wire [2:0] widget_auto_in_a_bits_opcode;
	wire [2:0] widget_auto_in_a_bits_param;
	wire [3:0] widget_auto_in_a_bits_size;
	wire [1:0] widget_auto_in_a_bits_source;
	wire [31:0] widget_auto_in_a_bits_address;
	wire [3:0] widget_auto_in_a_bits_mask;
	wire [31:0] widget_auto_in_a_bits_data;
	wire widget_auto_in_a_bits_corrupt;
	wire widget_auto_in_d_ready;
	wire widget_auto_in_d_valid;
	wire [2:0] widget_auto_in_d_bits_opcode;
	wire [1:0] widget_auto_in_d_bits_param;
	wire [3:0] widget_auto_in_d_bits_size;
	wire [1:0] widget_auto_in_d_bits_source;
	wire widget_auto_in_d_bits_sink;
	wire widget_auto_in_d_bits_denied;
	wire [31:0] widget_auto_in_d_bits_data;
	wire widget_auto_in_d_bits_corrupt;
	wire widget_auto_out_a_ready;
	wire widget_auto_out_a_valid;
	wire [2:0] widget_auto_out_a_bits_opcode;
	wire [2:0] widget_auto_out_a_bits_param;
	wire [3:0] widget_auto_out_a_bits_size;
	wire [1:0] widget_auto_out_a_bits_source;
	wire [31:0] widget_auto_out_a_bits_address;
	wire [3:0] widget_auto_out_a_bits_mask;
	wire [31:0] widget_auto_out_a_bits_data;
	wire widget_auto_out_a_bits_corrupt;
	wire widget_auto_out_d_ready;
	wire widget_auto_out_d_valid;
	wire [2:0] widget_auto_out_d_bits_opcode;
	wire [1:0] widget_auto_out_d_bits_param;
	wire [3:0] widget_auto_out_d_bits_size;
	wire [1:0] widget_auto_out_d_bits_source;
	wire widget_auto_out_d_bits_sink;
	wire widget_auto_out_d_bits_denied;
	wire [31:0] widget_auto_out_d_bits_data;
	wire widget_auto_out_d_bits_corrupt;
	TLWidthWidget widget(
		.auto_in_a_ready(widget_auto_in_a_ready),
		.auto_in_a_valid(widget_auto_in_a_valid),
		.auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(widget_auto_in_a_bits_param),
		.auto_in_a_bits_size(widget_auto_in_a_bits_size),
		.auto_in_a_bits_source(widget_auto_in_a_bits_source),
		.auto_in_a_bits_address(widget_auto_in_a_bits_address),
		.auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
		.auto_in_a_bits_data(widget_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(widget_auto_in_a_bits_corrupt),
		.auto_in_d_ready(widget_auto_in_d_ready),
		.auto_in_d_valid(widget_auto_in_d_valid),
		.auto_in_d_bits_opcode(widget_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(widget_auto_in_d_bits_param),
		.auto_in_d_bits_size(widget_auto_in_d_bits_size),
		.auto_in_d_bits_source(widget_auto_in_d_bits_source),
		.auto_in_d_bits_sink(widget_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(widget_auto_in_d_bits_denied),
		.auto_in_d_bits_data(widget_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(widget_auto_in_d_bits_corrupt),
		.auto_out_a_ready(widget_auto_out_a_ready),
		.auto_out_a_valid(widget_auto_out_a_valid),
		.auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(widget_auto_out_a_bits_param),
		.auto_out_a_bits_size(widget_auto_out_a_bits_size),
		.auto_out_a_bits_source(widget_auto_out_a_bits_source),
		.auto_out_a_bits_address(widget_auto_out_a_bits_address),
		.auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
		.auto_out_a_bits_data(widget_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(widget_auto_out_a_bits_corrupt),
		.auto_out_d_ready(widget_auto_out_d_ready),
		.auto_out_d_valid(widget_auto_out_d_valid),
		.auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(widget_auto_out_d_bits_param),
		.auto_out_d_bits_size(widget_auto_out_d_bits_size),
		.auto_out_d_bits_source(widget_auto_out_d_bits_source),
		.auto_out_d_bits_sink(widget_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(widget_auto_out_d_bits_denied),
		.auto_out_d_bits_data(widget_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(widget_auto_out_d_bits_corrupt)
	);
	assign auto_widget_in_a_ready = widget_auto_in_a_ready;
	assign auto_widget_in_d_valid = widget_auto_in_d_valid;
	assign auto_widget_in_d_bits_opcode = widget_auto_in_d_bits_opcode;
	assign auto_widget_in_d_bits_param = widget_auto_in_d_bits_param;
	assign auto_widget_in_d_bits_size = widget_auto_in_d_bits_size;
	assign auto_widget_in_d_bits_source = widget_auto_in_d_bits_source;
	assign auto_widget_in_d_bits_sink = widget_auto_in_d_bits_sink;
	assign auto_widget_in_d_bits_denied = widget_auto_in_d_bits_denied;
	assign auto_widget_in_d_bits_data = widget_auto_in_d_bits_data;
	assign auto_widget_in_d_bits_corrupt = widget_auto_in_d_bits_corrupt;
	assign auto_bus_xing_out_a_valid = widget_auto_out_a_valid;
	assign auto_bus_xing_out_a_bits_opcode = widget_auto_out_a_bits_opcode;
	assign auto_bus_xing_out_a_bits_param = widget_auto_out_a_bits_param;
	assign auto_bus_xing_out_a_bits_size = widget_auto_out_a_bits_size;
	assign auto_bus_xing_out_a_bits_source = widget_auto_out_a_bits_source;
	assign auto_bus_xing_out_a_bits_address = widget_auto_out_a_bits_address;
	assign auto_bus_xing_out_a_bits_mask = widget_auto_out_a_bits_mask;
	assign auto_bus_xing_out_a_bits_data = widget_auto_out_a_bits_data;
	assign auto_bus_xing_out_a_bits_corrupt = widget_auto_out_a_bits_corrupt;
	assign auto_bus_xing_out_d_ready = widget_auto_out_d_ready;
	assign widget_auto_in_a_valid = auto_widget_in_a_valid;
	assign widget_auto_in_a_bits_opcode = auto_widget_in_a_bits_opcode;
	assign widget_auto_in_a_bits_param = auto_widget_in_a_bits_param;
	assign widget_auto_in_a_bits_size = auto_widget_in_a_bits_size;
	assign widget_auto_in_a_bits_source = auto_widget_in_a_bits_source;
	assign widget_auto_in_a_bits_address = auto_widget_in_a_bits_address;
	assign widget_auto_in_a_bits_mask = auto_widget_in_a_bits_mask;
	assign widget_auto_in_a_bits_data = auto_widget_in_a_bits_data;
	assign widget_auto_in_a_bits_corrupt = auto_widget_in_a_bits_corrupt;
	assign widget_auto_in_d_ready = auto_widget_in_d_ready;
	assign widget_auto_out_a_ready = auto_bus_xing_out_a_ready;
	assign widget_auto_out_d_valid = auto_bus_xing_out_d_valid;
	assign widget_auto_out_d_bits_opcode = auto_bus_xing_out_d_bits_opcode;
	assign widget_auto_out_d_bits_param = auto_bus_xing_out_d_bits_param;
	assign widget_auto_out_d_bits_size = auto_bus_xing_out_d_bits_size;
	assign widget_auto_out_d_bits_source = auto_bus_xing_out_d_bits_source;
	assign widget_auto_out_d_bits_sink = auto_bus_xing_out_d_bits_sink;
	assign widget_auto_out_d_bits_denied = auto_bus_xing_out_d_bits_denied;
	assign widget_auto_out_d_bits_data = auto_bus_xing_out_d_bits_data;
	assign widget_auto_out_d_bits_corrupt = auto_bus_xing_out_d_bits_corrupt;
endmodule
module TLWidthWidget_1 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module TLInterconnectCoupler_1 (
	auto_widget_out_a_ready,
	auto_widget_out_a_valid,
	auto_widget_out_a_bits_opcode,
	auto_widget_out_a_bits_param,
	auto_widget_out_a_bits_size,
	auto_widget_out_a_bits_source,
	auto_widget_out_a_bits_address,
	auto_widget_out_a_bits_mask,
	auto_widget_out_a_bits_data,
	auto_widget_out_a_bits_corrupt,
	auto_widget_out_d_ready,
	auto_widget_out_d_valid,
	auto_widget_out_d_bits_opcode,
	auto_widget_out_d_bits_param,
	auto_widget_out_d_bits_size,
	auto_widget_out_d_bits_sink,
	auto_widget_out_d_bits_denied,
	auto_widget_out_d_bits_data,
	auto_widget_out_d_bits_corrupt,
	auto_bus_xing_in_a_ready,
	auto_bus_xing_in_a_valid,
	auto_bus_xing_in_a_bits_opcode,
	auto_bus_xing_in_a_bits_param,
	auto_bus_xing_in_a_bits_size,
	auto_bus_xing_in_a_bits_source,
	auto_bus_xing_in_a_bits_address,
	auto_bus_xing_in_a_bits_mask,
	auto_bus_xing_in_a_bits_data,
	auto_bus_xing_in_a_bits_corrupt,
	auto_bus_xing_in_d_ready,
	auto_bus_xing_in_d_valid,
	auto_bus_xing_in_d_bits_opcode,
	auto_bus_xing_in_d_bits_param,
	auto_bus_xing_in_d_bits_size,
	auto_bus_xing_in_d_bits_sink,
	auto_bus_xing_in_d_bits_denied,
	auto_bus_xing_in_d_bits_data,
	auto_bus_xing_in_d_bits_corrupt
);
	input auto_widget_out_a_ready;
	output wire auto_widget_out_a_valid;
	output wire [2:0] auto_widget_out_a_bits_opcode;
	output wire [2:0] auto_widget_out_a_bits_param;
	output wire [3:0] auto_widget_out_a_bits_size;
	output wire auto_widget_out_a_bits_source;
	output wire [31:0] auto_widget_out_a_bits_address;
	output wire [3:0] auto_widget_out_a_bits_mask;
	output wire [31:0] auto_widget_out_a_bits_data;
	output wire auto_widget_out_a_bits_corrupt;
	output wire auto_widget_out_d_ready;
	input auto_widget_out_d_valid;
	input [2:0] auto_widget_out_d_bits_opcode;
	input [1:0] auto_widget_out_d_bits_param;
	input [3:0] auto_widget_out_d_bits_size;
	input auto_widget_out_d_bits_sink;
	input auto_widget_out_d_bits_denied;
	input [31:0] auto_widget_out_d_bits_data;
	input auto_widget_out_d_bits_corrupt;
	output wire auto_bus_xing_in_a_ready;
	input auto_bus_xing_in_a_valid;
	input [2:0] auto_bus_xing_in_a_bits_opcode;
	input [2:0] auto_bus_xing_in_a_bits_param;
	input [3:0] auto_bus_xing_in_a_bits_size;
	input auto_bus_xing_in_a_bits_source;
	input [31:0] auto_bus_xing_in_a_bits_address;
	input [3:0] auto_bus_xing_in_a_bits_mask;
	input [31:0] auto_bus_xing_in_a_bits_data;
	input auto_bus_xing_in_a_bits_corrupt;
	input auto_bus_xing_in_d_ready;
	output wire auto_bus_xing_in_d_valid;
	output wire [2:0] auto_bus_xing_in_d_bits_opcode;
	output wire [1:0] auto_bus_xing_in_d_bits_param;
	output wire [3:0] auto_bus_xing_in_d_bits_size;
	output wire auto_bus_xing_in_d_bits_sink;
	output wire auto_bus_xing_in_d_bits_denied;
	output wire [31:0] auto_bus_xing_in_d_bits_data;
	output wire auto_bus_xing_in_d_bits_corrupt;
	wire widget_auto_in_a_ready;
	wire widget_auto_in_a_valid;
	wire [2:0] widget_auto_in_a_bits_opcode;
	wire [2:0] widget_auto_in_a_bits_param;
	wire [3:0] widget_auto_in_a_bits_size;
	wire widget_auto_in_a_bits_source;
	wire [31:0] widget_auto_in_a_bits_address;
	wire [3:0] widget_auto_in_a_bits_mask;
	wire [31:0] widget_auto_in_a_bits_data;
	wire widget_auto_in_a_bits_corrupt;
	wire widget_auto_in_d_ready;
	wire widget_auto_in_d_valid;
	wire [2:0] widget_auto_in_d_bits_opcode;
	wire [1:0] widget_auto_in_d_bits_param;
	wire [3:0] widget_auto_in_d_bits_size;
	wire widget_auto_in_d_bits_sink;
	wire widget_auto_in_d_bits_denied;
	wire [31:0] widget_auto_in_d_bits_data;
	wire widget_auto_in_d_bits_corrupt;
	wire widget_auto_out_a_ready;
	wire widget_auto_out_a_valid;
	wire [2:0] widget_auto_out_a_bits_opcode;
	wire [2:0] widget_auto_out_a_bits_param;
	wire [3:0] widget_auto_out_a_bits_size;
	wire widget_auto_out_a_bits_source;
	wire [31:0] widget_auto_out_a_bits_address;
	wire [3:0] widget_auto_out_a_bits_mask;
	wire [31:0] widget_auto_out_a_bits_data;
	wire widget_auto_out_a_bits_corrupt;
	wire widget_auto_out_d_ready;
	wire widget_auto_out_d_valid;
	wire [2:0] widget_auto_out_d_bits_opcode;
	wire [1:0] widget_auto_out_d_bits_param;
	wire [3:0] widget_auto_out_d_bits_size;
	wire widget_auto_out_d_bits_sink;
	wire widget_auto_out_d_bits_denied;
	wire [31:0] widget_auto_out_d_bits_data;
	wire widget_auto_out_d_bits_corrupt;
	TLWidthWidget_1 widget(
		.auto_in_a_ready(widget_auto_in_a_ready),
		.auto_in_a_valid(widget_auto_in_a_valid),
		.auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(widget_auto_in_a_bits_param),
		.auto_in_a_bits_size(widget_auto_in_a_bits_size),
		.auto_in_a_bits_source(widget_auto_in_a_bits_source),
		.auto_in_a_bits_address(widget_auto_in_a_bits_address),
		.auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
		.auto_in_a_bits_data(widget_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(widget_auto_in_a_bits_corrupt),
		.auto_in_d_ready(widget_auto_in_d_ready),
		.auto_in_d_valid(widget_auto_in_d_valid),
		.auto_in_d_bits_opcode(widget_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(widget_auto_in_d_bits_param),
		.auto_in_d_bits_size(widget_auto_in_d_bits_size),
		.auto_in_d_bits_sink(widget_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(widget_auto_in_d_bits_denied),
		.auto_in_d_bits_data(widget_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(widget_auto_in_d_bits_corrupt),
		.auto_out_a_ready(widget_auto_out_a_ready),
		.auto_out_a_valid(widget_auto_out_a_valid),
		.auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(widget_auto_out_a_bits_param),
		.auto_out_a_bits_size(widget_auto_out_a_bits_size),
		.auto_out_a_bits_source(widget_auto_out_a_bits_source),
		.auto_out_a_bits_address(widget_auto_out_a_bits_address),
		.auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
		.auto_out_a_bits_data(widget_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(widget_auto_out_a_bits_corrupt),
		.auto_out_d_ready(widget_auto_out_d_ready),
		.auto_out_d_valid(widget_auto_out_d_valid),
		.auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(widget_auto_out_d_bits_param),
		.auto_out_d_bits_size(widget_auto_out_d_bits_size),
		.auto_out_d_bits_sink(widget_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(widget_auto_out_d_bits_denied),
		.auto_out_d_bits_data(widget_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(widget_auto_out_d_bits_corrupt)
	);
	assign auto_widget_out_a_valid = widget_auto_out_a_valid;
	assign auto_widget_out_a_bits_opcode = widget_auto_out_a_bits_opcode;
	assign auto_widget_out_a_bits_param = widget_auto_out_a_bits_param;
	assign auto_widget_out_a_bits_size = widget_auto_out_a_bits_size;
	assign auto_widget_out_a_bits_source = widget_auto_out_a_bits_source;
	assign auto_widget_out_a_bits_address = widget_auto_out_a_bits_address;
	assign auto_widget_out_a_bits_mask = widget_auto_out_a_bits_mask;
	assign auto_widget_out_a_bits_data = widget_auto_out_a_bits_data;
	assign auto_widget_out_a_bits_corrupt = widget_auto_out_a_bits_corrupt;
	assign auto_widget_out_d_ready = widget_auto_out_d_ready;
	assign auto_bus_xing_in_a_ready = widget_auto_in_a_ready;
	assign auto_bus_xing_in_d_valid = widget_auto_in_d_valid;
	assign auto_bus_xing_in_d_bits_opcode = widget_auto_in_d_bits_opcode;
	assign auto_bus_xing_in_d_bits_param = widget_auto_in_d_bits_param;
	assign auto_bus_xing_in_d_bits_size = widget_auto_in_d_bits_size;
	assign auto_bus_xing_in_d_bits_sink = widget_auto_in_d_bits_sink;
	assign auto_bus_xing_in_d_bits_denied = widget_auto_in_d_bits_denied;
	assign auto_bus_xing_in_d_bits_data = widget_auto_in_d_bits_data;
	assign auto_bus_xing_in_d_bits_corrupt = widget_auto_in_d_bits_corrupt;
	assign widget_auto_in_a_valid = auto_bus_xing_in_a_valid;
	assign widget_auto_in_a_bits_opcode = auto_bus_xing_in_a_bits_opcode;
	assign widget_auto_in_a_bits_param = auto_bus_xing_in_a_bits_param;
	assign widget_auto_in_a_bits_size = auto_bus_xing_in_a_bits_size;
	assign widget_auto_in_a_bits_source = auto_bus_xing_in_a_bits_source;
	assign widget_auto_in_a_bits_address = auto_bus_xing_in_a_bits_address;
	assign widget_auto_in_a_bits_mask = auto_bus_xing_in_a_bits_mask;
	assign widget_auto_in_a_bits_data = auto_bus_xing_in_a_bits_data;
	assign widget_auto_in_a_bits_corrupt = auto_bus_xing_in_a_bits_corrupt;
	assign widget_auto_in_d_ready = auto_bus_xing_in_d_ready;
	assign widget_auto_out_a_ready = auto_widget_out_a_ready;
	assign widget_auto_out_d_valid = auto_widget_out_d_valid;
	assign widget_auto_out_d_bits_opcode = auto_widget_out_d_bits_opcode;
	assign widget_auto_out_d_bits_param = auto_widget_out_d_bits_param;
	assign widget_auto_out_d_bits_size = auto_widget_out_d_bits_size;
	assign widget_auto_out_d_bits_sink = auto_widget_out_d_bits_sink;
	assign widget_auto_out_d_bits_denied = auto_widget_out_d_bits_denied;
	assign widget_auto_out_d_bits_data = auto_widget_out_d_bits_data;
	assign widget_auto_out_d_bits_corrupt = auto_widget_out_d_bits_corrupt;
endmodule
module TLInterconnectCoupler_2 (
	auto_tl_master_clock_xing_in_a_ready,
	auto_tl_master_clock_xing_in_a_valid,
	auto_tl_master_clock_xing_in_a_bits_opcode,
	auto_tl_master_clock_xing_in_a_bits_param,
	auto_tl_master_clock_xing_in_a_bits_size,
	auto_tl_master_clock_xing_in_a_bits_source,
	auto_tl_master_clock_xing_in_a_bits_address,
	auto_tl_master_clock_xing_in_a_bits_mask,
	auto_tl_master_clock_xing_in_a_bits_data,
	auto_tl_master_clock_xing_in_a_bits_corrupt,
	auto_tl_master_clock_xing_in_d_ready,
	auto_tl_master_clock_xing_in_d_valid,
	auto_tl_master_clock_xing_in_d_bits_opcode,
	auto_tl_master_clock_xing_in_d_bits_param,
	auto_tl_master_clock_xing_in_d_bits_size,
	auto_tl_master_clock_xing_in_d_bits_source,
	auto_tl_master_clock_xing_in_d_bits_sink,
	auto_tl_master_clock_xing_in_d_bits_denied,
	auto_tl_master_clock_xing_in_d_bits_data,
	auto_tl_master_clock_xing_in_d_bits_corrupt,
	auto_tl_out_a_ready,
	auto_tl_out_a_valid,
	auto_tl_out_a_bits_opcode,
	auto_tl_out_a_bits_param,
	auto_tl_out_a_bits_size,
	auto_tl_out_a_bits_source,
	auto_tl_out_a_bits_address,
	auto_tl_out_a_bits_mask,
	auto_tl_out_a_bits_data,
	auto_tl_out_a_bits_corrupt,
	auto_tl_out_d_ready,
	auto_tl_out_d_valid,
	auto_tl_out_d_bits_opcode,
	auto_tl_out_d_bits_param,
	auto_tl_out_d_bits_size,
	auto_tl_out_d_bits_source,
	auto_tl_out_d_bits_sink,
	auto_tl_out_d_bits_denied,
	auto_tl_out_d_bits_data,
	auto_tl_out_d_bits_corrupt
);
	output wire auto_tl_master_clock_xing_in_a_ready;
	input auto_tl_master_clock_xing_in_a_valid;
	input [2:0] auto_tl_master_clock_xing_in_a_bits_opcode;
	input [2:0] auto_tl_master_clock_xing_in_a_bits_param;
	input [3:0] auto_tl_master_clock_xing_in_a_bits_size;
	input auto_tl_master_clock_xing_in_a_bits_source;
	input [31:0] auto_tl_master_clock_xing_in_a_bits_address;
	input [3:0] auto_tl_master_clock_xing_in_a_bits_mask;
	input [31:0] auto_tl_master_clock_xing_in_a_bits_data;
	input auto_tl_master_clock_xing_in_a_bits_corrupt;
	input auto_tl_master_clock_xing_in_d_ready;
	output wire auto_tl_master_clock_xing_in_d_valid;
	output wire [2:0] auto_tl_master_clock_xing_in_d_bits_opcode;
	output wire [1:0] auto_tl_master_clock_xing_in_d_bits_param;
	output wire [3:0] auto_tl_master_clock_xing_in_d_bits_size;
	output wire auto_tl_master_clock_xing_in_d_bits_source;
	output wire auto_tl_master_clock_xing_in_d_bits_sink;
	output wire auto_tl_master_clock_xing_in_d_bits_denied;
	output wire [31:0] auto_tl_master_clock_xing_in_d_bits_data;
	output wire auto_tl_master_clock_xing_in_d_bits_corrupt;
	input auto_tl_out_a_ready;
	output wire auto_tl_out_a_valid;
	output wire [2:0] auto_tl_out_a_bits_opcode;
	output wire [2:0] auto_tl_out_a_bits_param;
	output wire [3:0] auto_tl_out_a_bits_size;
	output wire auto_tl_out_a_bits_source;
	output wire [31:0] auto_tl_out_a_bits_address;
	output wire [3:0] auto_tl_out_a_bits_mask;
	output wire [31:0] auto_tl_out_a_bits_data;
	output wire auto_tl_out_a_bits_corrupt;
	output wire auto_tl_out_d_ready;
	input auto_tl_out_d_valid;
	input [2:0] auto_tl_out_d_bits_opcode;
	input [1:0] auto_tl_out_d_bits_param;
	input [3:0] auto_tl_out_d_bits_size;
	input auto_tl_out_d_bits_source;
	input auto_tl_out_d_bits_sink;
	input auto_tl_out_d_bits_denied;
	input [31:0] auto_tl_out_d_bits_data;
	input auto_tl_out_d_bits_corrupt;
	assign auto_tl_master_clock_xing_in_a_ready = auto_tl_out_a_ready;
	assign auto_tl_master_clock_xing_in_d_valid = auto_tl_out_d_valid;
	assign auto_tl_master_clock_xing_in_d_bits_opcode = auto_tl_out_d_bits_opcode;
	assign auto_tl_master_clock_xing_in_d_bits_param = auto_tl_out_d_bits_param;
	assign auto_tl_master_clock_xing_in_d_bits_size = auto_tl_out_d_bits_size;
	assign auto_tl_master_clock_xing_in_d_bits_source = auto_tl_out_d_bits_source;
	assign auto_tl_master_clock_xing_in_d_bits_sink = auto_tl_out_d_bits_sink;
	assign auto_tl_master_clock_xing_in_d_bits_denied = auto_tl_out_d_bits_denied;
	assign auto_tl_master_clock_xing_in_d_bits_data = auto_tl_out_d_bits_data;
	assign auto_tl_master_clock_xing_in_d_bits_corrupt = auto_tl_out_d_bits_corrupt;
	assign auto_tl_out_a_valid = auto_tl_master_clock_xing_in_a_valid;
	assign auto_tl_out_a_bits_opcode = auto_tl_master_clock_xing_in_a_bits_opcode;
	assign auto_tl_out_a_bits_param = auto_tl_master_clock_xing_in_a_bits_param;
	assign auto_tl_out_a_bits_size = auto_tl_master_clock_xing_in_a_bits_size;
	assign auto_tl_out_a_bits_source = auto_tl_master_clock_xing_in_a_bits_source;
	assign auto_tl_out_a_bits_address = auto_tl_master_clock_xing_in_a_bits_address;
	assign auto_tl_out_a_bits_mask = auto_tl_master_clock_xing_in_a_bits_mask;
	assign auto_tl_out_a_bits_data = auto_tl_master_clock_xing_in_a_bits_data;
	assign auto_tl_out_a_bits_corrupt = auto_tl_master_clock_xing_in_a_bits_corrupt;
	assign auto_tl_out_d_ready = auto_tl_master_clock_xing_in_d_ready;
endmodule
module SystemBus (
	auto_coupler_from_tile_tl_master_clock_xing_in_a_ready,
	auto_coupler_from_tile_tl_master_clock_xing_in_a_valid,
	auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode,
	auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param,
	auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size,
	auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source,
	auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address,
	auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask,
	auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data,
	auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_corrupt,
	auto_coupler_from_tile_tl_master_clock_xing_in_d_ready,
	auto_coupler_from_tile_tl_master_clock_xing_in_d_valid,
	auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode,
	auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param,
	auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size,
	auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source,
	auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink,
	auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied,
	auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data,
	auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_corrupt,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data,
	auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data,
	auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt,
	auto_fixedClockNode_out_1_clock,
	auto_fixedClockNode_out_1_reset,
	auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock,
	auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset
);
	output wire auto_coupler_from_tile_tl_master_clock_xing_in_a_ready;
	input auto_coupler_from_tile_tl_master_clock_xing_in_a_valid;
	input [2:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode;
	input [2:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param;
	input [3:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size;
	input auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source;
	input [31:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address;
	input [3:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask;
	input [31:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data;
	input auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_corrupt;
	input auto_coupler_from_tile_tl_master_clock_xing_in_d_ready;
	output wire auto_coupler_from_tile_tl_master_clock_xing_in_d_valid;
	output wire [2:0] auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode;
	output wire [1:0] auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param;
	output wire [3:0] auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size;
	output wire auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source;
	output wire auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink;
	output wire auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied;
	output wire [31:0] auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data;
	output wire auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt;
	output wire auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready;
	input auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid;
	input [2:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode;
	input [2:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param;
	input [3:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size;
	input auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source;
	input [31:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address;
	input [3:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask;
	input [31:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data;
	input auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_corrupt;
	input auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready;
	output wire auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid;
	output wire [2:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode;
	output wire [1:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param;
	output wire [3:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size;
	output wire auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink;
	output wire auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied;
	output wire [31:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data;
	output wire auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt;
	input auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready;
	output wire auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid;
	output wire [2:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode;
	output wire [2:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param;
	output wire [3:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size;
	output wire [1:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source;
	output wire [31:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address;
	output wire [3:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask;
	output wire [31:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data;
	output wire auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt;
	output wire auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready;
	input auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid;
	input [2:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode;
	input [1:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param;
	input [3:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size;
	input [1:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source;
	input auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink;
	input auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied;
	input [31:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data;
	input auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt;
	output wire auto_fixedClockNode_out_1_clock;
	output wire auto_fixedClockNode_out_1_reset;
	input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock;
	input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset;
	wire subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_clock;
	wire subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_reset;
	wire subsystem_sbus_clock_groups_auto_out_member_subsystem_sbus_0_clock;
	wire subsystem_sbus_clock_groups_auto_out_member_subsystem_sbus_0_reset;
	wire clockGroup_auto_in_member_subsystem_sbus_0_clock;
	wire clockGroup_auto_in_member_subsystem_sbus_0_reset;
	wire clockGroup_auto_out_clock;
	wire clockGroup_auto_out_reset;
	wire fixedClockNode_auto_in_clock;
	wire fixedClockNode_auto_in_reset;
	wire fixedClockNode_auto_out_2_clock;
	wire fixedClockNode_auto_out_2_reset;
	wire fixedClockNode_auto_out_0_clock;
	wire fixedClockNode_auto_out_0_reset;
	wire system_bus_xbar_clock;
	wire system_bus_xbar_reset;
	wire system_bus_xbar_auto_in_1_a_ready;
	wire system_bus_xbar_auto_in_1_a_valid;
	wire [2:0] system_bus_xbar_auto_in_1_a_bits_opcode;
	wire [2:0] system_bus_xbar_auto_in_1_a_bits_param;
	wire [3:0] system_bus_xbar_auto_in_1_a_bits_size;
	wire system_bus_xbar_auto_in_1_a_bits_source;
	wire [31:0] system_bus_xbar_auto_in_1_a_bits_address;
	wire [3:0] system_bus_xbar_auto_in_1_a_bits_mask;
	wire [31:0] system_bus_xbar_auto_in_1_a_bits_data;
	wire system_bus_xbar_auto_in_1_a_bits_corrupt;
	wire system_bus_xbar_auto_in_1_d_ready;
	wire system_bus_xbar_auto_in_1_d_valid;
	wire [2:0] system_bus_xbar_auto_in_1_d_bits_opcode;
	wire [1:0] system_bus_xbar_auto_in_1_d_bits_param;
	wire [3:0] system_bus_xbar_auto_in_1_d_bits_size;
	wire system_bus_xbar_auto_in_1_d_bits_source;
	wire system_bus_xbar_auto_in_1_d_bits_sink;
	wire system_bus_xbar_auto_in_1_d_bits_denied;
	wire [31:0] system_bus_xbar_auto_in_1_d_bits_data;
	wire system_bus_xbar_auto_in_1_d_bits_corrupt;
	wire system_bus_xbar_auto_in_0_a_ready;
	wire system_bus_xbar_auto_in_0_a_valid;
	wire [2:0] system_bus_xbar_auto_in_0_a_bits_opcode;
	wire [2:0] system_bus_xbar_auto_in_0_a_bits_param;
	wire [3:0] system_bus_xbar_auto_in_0_a_bits_size;
	wire system_bus_xbar_auto_in_0_a_bits_source;
	wire [31:0] system_bus_xbar_auto_in_0_a_bits_address;
	wire [3:0] system_bus_xbar_auto_in_0_a_bits_mask;
	wire [31:0] system_bus_xbar_auto_in_0_a_bits_data;
	wire system_bus_xbar_auto_in_0_a_bits_corrupt;
	wire system_bus_xbar_auto_in_0_d_ready;
	wire system_bus_xbar_auto_in_0_d_valid;
	wire [2:0] system_bus_xbar_auto_in_0_d_bits_opcode;
	wire [1:0] system_bus_xbar_auto_in_0_d_bits_param;
	wire [3:0] system_bus_xbar_auto_in_0_d_bits_size;
	wire system_bus_xbar_auto_in_0_d_bits_sink;
	wire system_bus_xbar_auto_in_0_d_bits_denied;
	wire [31:0] system_bus_xbar_auto_in_0_d_bits_data;
	wire system_bus_xbar_auto_in_0_d_bits_corrupt;
	wire system_bus_xbar_auto_out_a_ready;
	wire system_bus_xbar_auto_out_a_valid;
	wire [2:0] system_bus_xbar_auto_out_a_bits_opcode;
	wire [2:0] system_bus_xbar_auto_out_a_bits_param;
	wire [3:0] system_bus_xbar_auto_out_a_bits_size;
	wire [1:0] system_bus_xbar_auto_out_a_bits_source;
	wire [31:0] system_bus_xbar_auto_out_a_bits_address;
	wire [3:0] system_bus_xbar_auto_out_a_bits_mask;
	wire [31:0] system_bus_xbar_auto_out_a_bits_data;
	wire system_bus_xbar_auto_out_a_bits_corrupt;
	wire system_bus_xbar_auto_out_d_ready;
	wire system_bus_xbar_auto_out_d_valid;
	wire [2:0] system_bus_xbar_auto_out_d_bits_opcode;
	wire [1:0] system_bus_xbar_auto_out_d_bits_param;
	wire [3:0] system_bus_xbar_auto_out_d_bits_size;
	wire [1:0] system_bus_xbar_auto_out_d_bits_source;
	wire system_bus_xbar_auto_out_d_bits_sink;
	wire system_bus_xbar_auto_out_d_bits_denied;
	wire [31:0] system_bus_xbar_auto_out_d_bits_data;
	wire system_bus_xbar_auto_out_d_bits_corrupt;
	wire fixer_clock;
	wire fixer_reset;
	wire fixer_auto_in_1_a_ready;
	wire fixer_auto_in_1_a_valid;
	wire [2:0] fixer_auto_in_1_a_bits_opcode;
	wire [2:0] fixer_auto_in_1_a_bits_param;
	wire [3:0] fixer_auto_in_1_a_bits_size;
	wire fixer_auto_in_1_a_bits_source;
	wire [31:0] fixer_auto_in_1_a_bits_address;
	wire [3:0] fixer_auto_in_1_a_bits_mask;
	wire [31:0] fixer_auto_in_1_a_bits_data;
	wire fixer_auto_in_1_a_bits_corrupt;
	wire fixer_auto_in_1_d_ready;
	wire fixer_auto_in_1_d_valid;
	wire [2:0] fixer_auto_in_1_d_bits_opcode;
	wire [1:0] fixer_auto_in_1_d_bits_param;
	wire [3:0] fixer_auto_in_1_d_bits_size;
	wire fixer_auto_in_1_d_bits_source;
	wire fixer_auto_in_1_d_bits_sink;
	wire fixer_auto_in_1_d_bits_denied;
	wire [31:0] fixer_auto_in_1_d_bits_data;
	wire fixer_auto_in_1_d_bits_corrupt;
	wire fixer_auto_in_0_a_ready;
	wire fixer_auto_in_0_a_valid;
	wire [2:0] fixer_auto_in_0_a_bits_opcode;
	wire [2:0] fixer_auto_in_0_a_bits_param;
	wire [3:0] fixer_auto_in_0_a_bits_size;
	wire fixer_auto_in_0_a_bits_source;
	wire [31:0] fixer_auto_in_0_a_bits_address;
	wire [3:0] fixer_auto_in_0_a_bits_mask;
	wire [31:0] fixer_auto_in_0_a_bits_data;
	wire fixer_auto_in_0_a_bits_corrupt;
	wire fixer_auto_in_0_d_ready;
	wire fixer_auto_in_0_d_valid;
	wire [2:0] fixer_auto_in_0_d_bits_opcode;
	wire [1:0] fixer_auto_in_0_d_bits_param;
	wire [3:0] fixer_auto_in_0_d_bits_size;
	wire fixer_auto_in_0_d_bits_sink;
	wire fixer_auto_in_0_d_bits_denied;
	wire [31:0] fixer_auto_in_0_d_bits_data;
	wire fixer_auto_in_0_d_bits_corrupt;
	wire fixer_auto_out_1_a_ready;
	wire fixer_auto_out_1_a_valid;
	wire [2:0] fixer_auto_out_1_a_bits_opcode;
	wire [2:0] fixer_auto_out_1_a_bits_param;
	wire [3:0] fixer_auto_out_1_a_bits_size;
	wire fixer_auto_out_1_a_bits_source;
	wire [31:0] fixer_auto_out_1_a_bits_address;
	wire [3:0] fixer_auto_out_1_a_bits_mask;
	wire [31:0] fixer_auto_out_1_a_bits_data;
	wire fixer_auto_out_1_a_bits_corrupt;
	wire fixer_auto_out_1_d_ready;
	wire fixer_auto_out_1_d_valid;
	wire [2:0] fixer_auto_out_1_d_bits_opcode;
	wire [1:0] fixer_auto_out_1_d_bits_param;
	wire [3:0] fixer_auto_out_1_d_bits_size;
	wire fixer_auto_out_1_d_bits_source;
	wire fixer_auto_out_1_d_bits_sink;
	wire fixer_auto_out_1_d_bits_denied;
	wire [31:0] fixer_auto_out_1_d_bits_data;
	wire fixer_auto_out_1_d_bits_corrupt;
	wire fixer_auto_out_0_a_ready;
	wire fixer_auto_out_0_a_valid;
	wire [2:0] fixer_auto_out_0_a_bits_opcode;
	wire [2:0] fixer_auto_out_0_a_bits_param;
	wire [3:0] fixer_auto_out_0_a_bits_size;
	wire fixer_auto_out_0_a_bits_source;
	wire [31:0] fixer_auto_out_0_a_bits_address;
	wire [3:0] fixer_auto_out_0_a_bits_mask;
	wire [31:0] fixer_auto_out_0_a_bits_data;
	wire fixer_auto_out_0_a_bits_corrupt;
	wire fixer_auto_out_0_d_ready;
	wire fixer_auto_out_0_d_valid;
	wire [2:0] fixer_auto_out_0_d_bits_opcode;
	wire [1:0] fixer_auto_out_0_d_bits_param;
	wire [3:0] fixer_auto_out_0_d_bits_size;
	wire fixer_auto_out_0_d_bits_sink;
	wire fixer_auto_out_0_d_bits_denied;
	wire [31:0] fixer_auto_out_0_d_bits_data;
	wire fixer_auto_out_0_d_bits_corrupt;
	wire coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_ready;
	wire coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_valid;
	wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_opcode;
	wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_param;
	wire [3:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_size;
	wire [1:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_source;
	wire [31:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_address;
	wire [3:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_mask;
	wire [31:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_data;
	wire coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_corrupt;
	wire coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_ready;
	wire coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_valid;
	wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_opcode;
	wire [1:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_param;
	wire [3:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_size;
	wire [1:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_source;
	wire coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_sink;
	wire coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_denied;
	wire [31:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_data;
	wire coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_corrupt;
	wire coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_ready;
	wire coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_valid;
	wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_opcode;
	wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_param;
	wire [3:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_size;
	wire [1:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_source;
	wire [31:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_address;
	wire [3:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_mask;
	wire [31:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_data;
	wire coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_corrupt;
	wire coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_ready;
	wire coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_valid;
	wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_opcode;
	wire [1:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_param;
	wire [3:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_size;
	wire [1:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_source;
	wire coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_sink;
	wire coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_denied;
	wire [31:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_data;
	wire coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_corrupt;
	wire coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_ready;
	wire coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_valid;
	wire [2:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_opcode;
	wire [2:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_param;
	wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_size;
	wire coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_source;
	wire [31:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_address;
	wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_mask;
	wire [31:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_data;
	wire coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_corrupt;
	wire coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_ready;
	wire coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_valid;
	wire [2:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_opcode;
	wire [1:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_param;
	wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_size;
	wire coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_sink;
	wire coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_denied;
	wire [31:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_data;
	wire coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_corrupt;
	wire coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_ready;
	wire coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_valid;
	wire [2:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_opcode;
	wire [2:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_param;
	wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_size;
	wire coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_source;
	wire [31:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_address;
	wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_mask;
	wire [31:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_data;
	wire coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_corrupt;
	wire coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_ready;
	wire coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_valid;
	wire [2:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_opcode;
	wire [1:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_param;
	wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_size;
	wire coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_sink;
	wire coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_denied;
	wire [31:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_data;
	wire coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_corrupt;
	wire coupler_from_tile_auto_tl_master_clock_xing_in_a_ready;
	wire coupler_from_tile_auto_tl_master_clock_xing_in_a_valid;
	wire [2:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_opcode;
	wire [2:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_param;
	wire [3:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_size;
	wire coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_source;
	wire [31:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_address;
	wire [3:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_mask;
	wire [31:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_data;
	wire coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_corrupt;
	wire coupler_from_tile_auto_tl_master_clock_xing_in_d_ready;
	wire coupler_from_tile_auto_tl_master_clock_xing_in_d_valid;
	wire [2:0] coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_opcode;
	wire [1:0] coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_param;
	wire [3:0] coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_size;
	wire coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_source;
	wire coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_sink;
	wire coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_denied;
	wire [31:0] coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_data;
	wire coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_corrupt;
	wire coupler_from_tile_auto_tl_out_a_ready;
	wire coupler_from_tile_auto_tl_out_a_valid;
	wire [2:0] coupler_from_tile_auto_tl_out_a_bits_opcode;
	wire [2:0] coupler_from_tile_auto_tl_out_a_bits_param;
	wire [3:0] coupler_from_tile_auto_tl_out_a_bits_size;
	wire coupler_from_tile_auto_tl_out_a_bits_source;
	wire [31:0] coupler_from_tile_auto_tl_out_a_bits_address;
	wire [3:0] coupler_from_tile_auto_tl_out_a_bits_mask;
	wire [31:0] coupler_from_tile_auto_tl_out_a_bits_data;
	wire coupler_from_tile_auto_tl_out_a_bits_corrupt;
	wire coupler_from_tile_auto_tl_out_d_ready;
	wire coupler_from_tile_auto_tl_out_d_valid;
	wire [2:0] coupler_from_tile_auto_tl_out_d_bits_opcode;
	wire [1:0] coupler_from_tile_auto_tl_out_d_bits_param;
	wire [3:0] coupler_from_tile_auto_tl_out_d_bits_size;
	wire coupler_from_tile_auto_tl_out_d_bits_source;
	wire coupler_from_tile_auto_tl_out_d_bits_sink;
	wire coupler_from_tile_auto_tl_out_d_bits_denied;
	wire [31:0] coupler_from_tile_auto_tl_out_d_bits_data;
	wire coupler_from_tile_auto_tl_out_d_bits_corrupt;
	ClockGroupAggregator subsystem_sbus_clock_groups(
		.auto_in_member_subsystem_sbus_0_clock(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_clock),
		.auto_in_member_subsystem_sbus_0_reset(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_reset),
		.auto_out_member_subsystem_sbus_0_clock(subsystem_sbus_clock_groups_auto_out_member_subsystem_sbus_0_clock),
		.auto_out_member_subsystem_sbus_0_reset(subsystem_sbus_clock_groups_auto_out_member_subsystem_sbus_0_reset)
	);
	ClockGroup clockGroup(
		.auto_in_member_subsystem_sbus_0_clock(clockGroup_auto_in_member_subsystem_sbus_0_clock),
		.auto_in_member_subsystem_sbus_0_reset(clockGroup_auto_in_member_subsystem_sbus_0_reset),
		.auto_out_clock(clockGroup_auto_out_clock),
		.auto_out_reset(clockGroup_auto_out_reset)
	);
	FixedClockBroadcast fixedClockNode(
		.auto_in_clock(fixedClockNode_auto_in_clock),
		.auto_in_reset(fixedClockNode_auto_in_reset),
		.auto_out_2_clock(fixedClockNode_auto_out_2_clock),
		.auto_out_2_reset(fixedClockNode_auto_out_2_reset),
		.auto_out_0_clock(fixedClockNode_auto_out_0_clock),
		.auto_out_0_reset(fixedClockNode_auto_out_0_reset)
	);
	TLXbar system_bus_xbar(
		.clock(system_bus_xbar_clock),
		.reset(system_bus_xbar_reset),
		.auto_in_1_a_ready(system_bus_xbar_auto_in_1_a_ready),
		.auto_in_1_a_valid(system_bus_xbar_auto_in_1_a_valid),
		.auto_in_1_a_bits_opcode(system_bus_xbar_auto_in_1_a_bits_opcode),
		.auto_in_1_a_bits_param(system_bus_xbar_auto_in_1_a_bits_param),
		.auto_in_1_a_bits_size(system_bus_xbar_auto_in_1_a_bits_size),
		.auto_in_1_a_bits_source(system_bus_xbar_auto_in_1_a_bits_source),
		.auto_in_1_a_bits_address(system_bus_xbar_auto_in_1_a_bits_address),
		.auto_in_1_a_bits_mask(system_bus_xbar_auto_in_1_a_bits_mask),
		.auto_in_1_a_bits_data(system_bus_xbar_auto_in_1_a_bits_data),
		.auto_in_1_a_bits_corrupt(system_bus_xbar_auto_in_1_a_bits_corrupt),
		.auto_in_1_d_ready(system_bus_xbar_auto_in_1_d_ready),
		.auto_in_1_d_valid(system_bus_xbar_auto_in_1_d_valid),
		.auto_in_1_d_bits_opcode(system_bus_xbar_auto_in_1_d_bits_opcode),
		.auto_in_1_d_bits_param(system_bus_xbar_auto_in_1_d_bits_param),
		.auto_in_1_d_bits_size(system_bus_xbar_auto_in_1_d_bits_size),
		.auto_in_1_d_bits_source(system_bus_xbar_auto_in_1_d_bits_source),
		.auto_in_1_d_bits_sink(system_bus_xbar_auto_in_1_d_bits_sink),
		.auto_in_1_d_bits_denied(system_bus_xbar_auto_in_1_d_bits_denied),
		.auto_in_1_d_bits_data(system_bus_xbar_auto_in_1_d_bits_data),
		.auto_in_1_d_bits_corrupt(system_bus_xbar_auto_in_1_d_bits_corrupt),
		.auto_in_0_a_ready(system_bus_xbar_auto_in_0_a_ready),
		.auto_in_0_a_valid(system_bus_xbar_auto_in_0_a_valid),
		.auto_in_0_a_bits_opcode(system_bus_xbar_auto_in_0_a_bits_opcode),
		.auto_in_0_a_bits_param(system_bus_xbar_auto_in_0_a_bits_param),
		.auto_in_0_a_bits_size(system_bus_xbar_auto_in_0_a_bits_size),
		.auto_in_0_a_bits_source(system_bus_xbar_auto_in_0_a_bits_source),
		.auto_in_0_a_bits_address(system_bus_xbar_auto_in_0_a_bits_address),
		.auto_in_0_a_bits_mask(system_bus_xbar_auto_in_0_a_bits_mask),
		.auto_in_0_a_bits_data(system_bus_xbar_auto_in_0_a_bits_data),
		.auto_in_0_a_bits_corrupt(system_bus_xbar_auto_in_0_a_bits_corrupt),
		.auto_in_0_d_ready(system_bus_xbar_auto_in_0_d_ready),
		.auto_in_0_d_valid(system_bus_xbar_auto_in_0_d_valid),
		.auto_in_0_d_bits_opcode(system_bus_xbar_auto_in_0_d_bits_opcode),
		.auto_in_0_d_bits_param(system_bus_xbar_auto_in_0_d_bits_param),
		.auto_in_0_d_bits_size(system_bus_xbar_auto_in_0_d_bits_size),
		.auto_in_0_d_bits_sink(system_bus_xbar_auto_in_0_d_bits_sink),
		.auto_in_0_d_bits_denied(system_bus_xbar_auto_in_0_d_bits_denied),
		.auto_in_0_d_bits_data(system_bus_xbar_auto_in_0_d_bits_data),
		.auto_in_0_d_bits_corrupt(system_bus_xbar_auto_in_0_d_bits_corrupt),
		.auto_out_a_ready(system_bus_xbar_auto_out_a_ready),
		.auto_out_a_valid(system_bus_xbar_auto_out_a_valid),
		.auto_out_a_bits_opcode(system_bus_xbar_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(system_bus_xbar_auto_out_a_bits_param),
		.auto_out_a_bits_size(system_bus_xbar_auto_out_a_bits_size),
		.auto_out_a_bits_source(system_bus_xbar_auto_out_a_bits_source),
		.auto_out_a_bits_address(system_bus_xbar_auto_out_a_bits_address),
		.auto_out_a_bits_mask(system_bus_xbar_auto_out_a_bits_mask),
		.auto_out_a_bits_data(system_bus_xbar_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(system_bus_xbar_auto_out_a_bits_corrupt),
		.auto_out_d_ready(system_bus_xbar_auto_out_d_ready),
		.auto_out_d_valid(system_bus_xbar_auto_out_d_valid),
		.auto_out_d_bits_opcode(system_bus_xbar_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(system_bus_xbar_auto_out_d_bits_param),
		.auto_out_d_bits_size(system_bus_xbar_auto_out_d_bits_size),
		.auto_out_d_bits_source(system_bus_xbar_auto_out_d_bits_source),
		.auto_out_d_bits_sink(system_bus_xbar_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(system_bus_xbar_auto_out_d_bits_denied),
		.auto_out_d_bits_data(system_bus_xbar_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(system_bus_xbar_auto_out_d_bits_corrupt)
	);
	TLFIFOFixer fixer(
		.clock(fixer_clock),
		.reset(fixer_reset),
		.auto_in_1_a_ready(fixer_auto_in_1_a_ready),
		.auto_in_1_a_valid(fixer_auto_in_1_a_valid),
		.auto_in_1_a_bits_opcode(fixer_auto_in_1_a_bits_opcode),
		.auto_in_1_a_bits_param(fixer_auto_in_1_a_bits_param),
		.auto_in_1_a_bits_size(fixer_auto_in_1_a_bits_size),
		.auto_in_1_a_bits_source(fixer_auto_in_1_a_bits_source),
		.auto_in_1_a_bits_address(fixer_auto_in_1_a_bits_address),
		.auto_in_1_a_bits_mask(fixer_auto_in_1_a_bits_mask),
		.auto_in_1_a_bits_data(fixer_auto_in_1_a_bits_data),
		.auto_in_1_a_bits_corrupt(fixer_auto_in_1_a_bits_corrupt),
		.auto_in_1_d_ready(fixer_auto_in_1_d_ready),
		.auto_in_1_d_valid(fixer_auto_in_1_d_valid),
		.auto_in_1_d_bits_opcode(fixer_auto_in_1_d_bits_opcode),
		.auto_in_1_d_bits_param(fixer_auto_in_1_d_bits_param),
		.auto_in_1_d_bits_size(fixer_auto_in_1_d_bits_size),
		.auto_in_1_d_bits_source(fixer_auto_in_1_d_bits_source),
		.auto_in_1_d_bits_sink(fixer_auto_in_1_d_bits_sink),
		.auto_in_1_d_bits_denied(fixer_auto_in_1_d_bits_denied),
		.auto_in_1_d_bits_data(fixer_auto_in_1_d_bits_data),
		.auto_in_1_d_bits_corrupt(fixer_auto_in_1_d_bits_corrupt),
		.auto_in_0_a_ready(fixer_auto_in_0_a_ready),
		.auto_in_0_a_valid(fixer_auto_in_0_a_valid),
		.auto_in_0_a_bits_opcode(fixer_auto_in_0_a_bits_opcode),
		.auto_in_0_a_bits_param(fixer_auto_in_0_a_bits_param),
		.auto_in_0_a_bits_size(fixer_auto_in_0_a_bits_size),
		.auto_in_0_a_bits_source(fixer_auto_in_0_a_bits_source),
		.auto_in_0_a_bits_address(fixer_auto_in_0_a_bits_address),
		.auto_in_0_a_bits_mask(fixer_auto_in_0_a_bits_mask),
		.auto_in_0_a_bits_data(fixer_auto_in_0_a_bits_data),
		.auto_in_0_a_bits_corrupt(fixer_auto_in_0_a_bits_corrupt),
		.auto_in_0_d_ready(fixer_auto_in_0_d_ready),
		.auto_in_0_d_valid(fixer_auto_in_0_d_valid),
		.auto_in_0_d_bits_opcode(fixer_auto_in_0_d_bits_opcode),
		.auto_in_0_d_bits_param(fixer_auto_in_0_d_bits_param),
		.auto_in_0_d_bits_size(fixer_auto_in_0_d_bits_size),
		.auto_in_0_d_bits_sink(fixer_auto_in_0_d_bits_sink),
		.auto_in_0_d_bits_denied(fixer_auto_in_0_d_bits_denied),
		.auto_in_0_d_bits_data(fixer_auto_in_0_d_bits_data),
		.auto_in_0_d_bits_corrupt(fixer_auto_in_0_d_bits_corrupt),
		.auto_out_1_a_ready(fixer_auto_out_1_a_ready),
		.auto_out_1_a_valid(fixer_auto_out_1_a_valid),
		.auto_out_1_a_bits_opcode(fixer_auto_out_1_a_bits_opcode),
		.auto_out_1_a_bits_param(fixer_auto_out_1_a_bits_param),
		.auto_out_1_a_bits_size(fixer_auto_out_1_a_bits_size),
		.auto_out_1_a_bits_source(fixer_auto_out_1_a_bits_source),
		.auto_out_1_a_bits_address(fixer_auto_out_1_a_bits_address),
		.auto_out_1_a_bits_mask(fixer_auto_out_1_a_bits_mask),
		.auto_out_1_a_bits_data(fixer_auto_out_1_a_bits_data),
		.auto_out_1_a_bits_corrupt(fixer_auto_out_1_a_bits_corrupt),
		.auto_out_1_d_ready(fixer_auto_out_1_d_ready),
		.auto_out_1_d_valid(fixer_auto_out_1_d_valid),
		.auto_out_1_d_bits_opcode(fixer_auto_out_1_d_bits_opcode),
		.auto_out_1_d_bits_param(fixer_auto_out_1_d_bits_param),
		.auto_out_1_d_bits_size(fixer_auto_out_1_d_bits_size),
		.auto_out_1_d_bits_source(fixer_auto_out_1_d_bits_source),
		.auto_out_1_d_bits_sink(fixer_auto_out_1_d_bits_sink),
		.auto_out_1_d_bits_denied(fixer_auto_out_1_d_bits_denied),
		.auto_out_1_d_bits_data(fixer_auto_out_1_d_bits_data),
		.auto_out_1_d_bits_corrupt(fixer_auto_out_1_d_bits_corrupt),
		.auto_out_0_a_ready(fixer_auto_out_0_a_ready),
		.auto_out_0_a_valid(fixer_auto_out_0_a_valid),
		.auto_out_0_a_bits_opcode(fixer_auto_out_0_a_bits_opcode),
		.auto_out_0_a_bits_param(fixer_auto_out_0_a_bits_param),
		.auto_out_0_a_bits_size(fixer_auto_out_0_a_bits_size),
		.auto_out_0_a_bits_source(fixer_auto_out_0_a_bits_source),
		.auto_out_0_a_bits_address(fixer_auto_out_0_a_bits_address),
		.auto_out_0_a_bits_mask(fixer_auto_out_0_a_bits_mask),
		.auto_out_0_a_bits_data(fixer_auto_out_0_a_bits_data),
		.auto_out_0_a_bits_corrupt(fixer_auto_out_0_a_bits_corrupt),
		.auto_out_0_d_ready(fixer_auto_out_0_d_ready),
		.auto_out_0_d_valid(fixer_auto_out_0_d_valid),
		.auto_out_0_d_bits_opcode(fixer_auto_out_0_d_bits_opcode),
		.auto_out_0_d_bits_param(fixer_auto_out_0_d_bits_param),
		.auto_out_0_d_bits_size(fixer_auto_out_0_d_bits_size),
		.auto_out_0_d_bits_sink(fixer_auto_out_0_d_bits_sink),
		.auto_out_0_d_bits_denied(fixer_auto_out_0_d_bits_denied),
		.auto_out_0_d_bits_data(fixer_auto_out_0_d_bits_data),
		.auto_out_0_d_bits_corrupt(fixer_auto_out_0_d_bits_corrupt)
	);
	TLInterconnectCoupler coupler_to_bus_named_subsystem_cbus(
		.auto_widget_in_a_ready(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_ready),
		.auto_widget_in_a_valid(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_valid),
		.auto_widget_in_a_bits_opcode(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_opcode),
		.auto_widget_in_a_bits_param(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_param),
		.auto_widget_in_a_bits_size(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_size),
		.auto_widget_in_a_bits_source(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_source),
		.auto_widget_in_a_bits_address(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_address),
		.auto_widget_in_a_bits_mask(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_mask),
		.auto_widget_in_a_bits_data(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_data),
		.auto_widget_in_a_bits_corrupt(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_corrupt),
		.auto_widget_in_d_ready(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_ready),
		.auto_widget_in_d_valid(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_valid),
		.auto_widget_in_d_bits_opcode(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_opcode),
		.auto_widget_in_d_bits_param(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_param),
		.auto_widget_in_d_bits_size(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_size),
		.auto_widget_in_d_bits_source(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_source),
		.auto_widget_in_d_bits_sink(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_sink),
		.auto_widget_in_d_bits_denied(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_denied),
		.auto_widget_in_d_bits_data(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_data),
		.auto_widget_in_d_bits_corrupt(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_corrupt),
		.auto_bus_xing_out_a_ready(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_ready),
		.auto_bus_xing_out_a_valid(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_valid),
		.auto_bus_xing_out_a_bits_opcode(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_opcode),
		.auto_bus_xing_out_a_bits_param(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_param),
		.auto_bus_xing_out_a_bits_size(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_size),
		.auto_bus_xing_out_a_bits_source(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_source),
		.auto_bus_xing_out_a_bits_address(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_address),
		.auto_bus_xing_out_a_bits_mask(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_mask),
		.auto_bus_xing_out_a_bits_data(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_data),
		.auto_bus_xing_out_a_bits_corrupt(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_corrupt),
		.auto_bus_xing_out_d_ready(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_ready),
		.auto_bus_xing_out_d_valid(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_valid),
		.auto_bus_xing_out_d_bits_opcode(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_opcode),
		.auto_bus_xing_out_d_bits_param(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_param),
		.auto_bus_xing_out_d_bits_size(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_size),
		.auto_bus_xing_out_d_bits_source(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_source),
		.auto_bus_xing_out_d_bits_sink(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_sink),
		.auto_bus_xing_out_d_bits_denied(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_denied),
		.auto_bus_xing_out_d_bits_data(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_data),
		.auto_bus_xing_out_d_bits_corrupt(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_corrupt)
	);
	TLInterconnectCoupler_1 coupler_from_bus_named_subsystem_fbus(
		.auto_widget_out_a_ready(coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_ready),
		.auto_widget_out_a_valid(coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_valid),
		.auto_widget_out_a_bits_opcode(coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_opcode),
		.auto_widget_out_a_bits_param(coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_param),
		.auto_widget_out_a_bits_size(coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_size),
		.auto_widget_out_a_bits_source(coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_source),
		.auto_widget_out_a_bits_address(coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_address),
		.auto_widget_out_a_bits_mask(coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_mask),
		.auto_widget_out_a_bits_data(coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_data),
		.auto_widget_out_a_bits_corrupt(coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_corrupt),
		.auto_widget_out_d_ready(coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_ready),
		.auto_widget_out_d_valid(coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_valid),
		.auto_widget_out_d_bits_opcode(coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_opcode),
		.auto_widget_out_d_bits_param(coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_param),
		.auto_widget_out_d_bits_size(coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_size),
		.auto_widget_out_d_bits_sink(coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_sink),
		.auto_widget_out_d_bits_denied(coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_denied),
		.auto_widget_out_d_bits_data(coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_data),
		.auto_widget_out_d_bits_corrupt(coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_corrupt),
		.auto_bus_xing_in_a_ready(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_ready),
		.auto_bus_xing_in_a_valid(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_valid),
		.auto_bus_xing_in_a_bits_opcode(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_opcode),
		.auto_bus_xing_in_a_bits_param(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_param),
		.auto_bus_xing_in_a_bits_size(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_size),
		.auto_bus_xing_in_a_bits_source(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_source),
		.auto_bus_xing_in_a_bits_address(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_address),
		.auto_bus_xing_in_a_bits_mask(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_mask),
		.auto_bus_xing_in_a_bits_data(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_data),
		.auto_bus_xing_in_a_bits_corrupt(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_corrupt),
		.auto_bus_xing_in_d_ready(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_ready),
		.auto_bus_xing_in_d_valid(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_valid),
		.auto_bus_xing_in_d_bits_opcode(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_opcode),
		.auto_bus_xing_in_d_bits_param(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_param),
		.auto_bus_xing_in_d_bits_size(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_size),
		.auto_bus_xing_in_d_bits_sink(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_sink),
		.auto_bus_xing_in_d_bits_denied(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_denied),
		.auto_bus_xing_in_d_bits_data(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_data),
		.auto_bus_xing_in_d_bits_corrupt(coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_corrupt)
	);
	TLInterconnectCoupler_2 coupler_from_tile(
		.auto_tl_master_clock_xing_in_a_ready(coupler_from_tile_auto_tl_master_clock_xing_in_a_ready),
		.auto_tl_master_clock_xing_in_a_valid(coupler_from_tile_auto_tl_master_clock_xing_in_a_valid),
		.auto_tl_master_clock_xing_in_a_bits_opcode(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_opcode),
		.auto_tl_master_clock_xing_in_a_bits_param(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_param),
		.auto_tl_master_clock_xing_in_a_bits_size(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_size),
		.auto_tl_master_clock_xing_in_a_bits_source(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_source),
		.auto_tl_master_clock_xing_in_a_bits_address(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_address),
		.auto_tl_master_clock_xing_in_a_bits_mask(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_mask),
		.auto_tl_master_clock_xing_in_a_bits_data(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_data),
		.auto_tl_master_clock_xing_in_a_bits_corrupt(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_corrupt),
		.auto_tl_master_clock_xing_in_d_ready(coupler_from_tile_auto_tl_master_clock_xing_in_d_ready),
		.auto_tl_master_clock_xing_in_d_valid(coupler_from_tile_auto_tl_master_clock_xing_in_d_valid),
		.auto_tl_master_clock_xing_in_d_bits_opcode(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_opcode),
		.auto_tl_master_clock_xing_in_d_bits_param(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_param),
		.auto_tl_master_clock_xing_in_d_bits_size(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_size),
		.auto_tl_master_clock_xing_in_d_bits_source(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_source),
		.auto_tl_master_clock_xing_in_d_bits_sink(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_sink),
		.auto_tl_master_clock_xing_in_d_bits_denied(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_denied),
		.auto_tl_master_clock_xing_in_d_bits_data(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_data),
		.auto_tl_master_clock_xing_in_d_bits_corrupt(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_corrupt),
		.auto_tl_out_a_ready(coupler_from_tile_auto_tl_out_a_ready),
		.auto_tl_out_a_valid(coupler_from_tile_auto_tl_out_a_valid),
		.auto_tl_out_a_bits_opcode(coupler_from_tile_auto_tl_out_a_bits_opcode),
		.auto_tl_out_a_bits_param(coupler_from_tile_auto_tl_out_a_bits_param),
		.auto_tl_out_a_bits_size(coupler_from_tile_auto_tl_out_a_bits_size),
		.auto_tl_out_a_bits_source(coupler_from_tile_auto_tl_out_a_bits_source),
		.auto_tl_out_a_bits_address(coupler_from_tile_auto_tl_out_a_bits_address),
		.auto_tl_out_a_bits_mask(coupler_from_tile_auto_tl_out_a_bits_mask),
		.auto_tl_out_a_bits_data(coupler_from_tile_auto_tl_out_a_bits_data),
		.auto_tl_out_a_bits_corrupt(coupler_from_tile_auto_tl_out_a_bits_corrupt),
		.auto_tl_out_d_ready(coupler_from_tile_auto_tl_out_d_ready),
		.auto_tl_out_d_valid(coupler_from_tile_auto_tl_out_d_valid),
		.auto_tl_out_d_bits_opcode(coupler_from_tile_auto_tl_out_d_bits_opcode),
		.auto_tl_out_d_bits_param(coupler_from_tile_auto_tl_out_d_bits_param),
		.auto_tl_out_d_bits_size(coupler_from_tile_auto_tl_out_d_bits_size),
		.auto_tl_out_d_bits_source(coupler_from_tile_auto_tl_out_d_bits_source),
		.auto_tl_out_d_bits_sink(coupler_from_tile_auto_tl_out_d_bits_sink),
		.auto_tl_out_d_bits_denied(coupler_from_tile_auto_tl_out_d_bits_denied),
		.auto_tl_out_d_bits_data(coupler_from_tile_auto_tl_out_d_bits_data),
		.auto_tl_out_d_bits_corrupt(coupler_from_tile_auto_tl_out_d_bits_corrupt)
	);
	assign auto_coupler_from_tile_tl_master_clock_xing_in_a_ready = coupler_from_tile_auto_tl_master_clock_xing_in_a_ready;
	assign auto_coupler_from_tile_tl_master_clock_xing_in_d_valid = coupler_from_tile_auto_tl_master_clock_xing_in_d_valid;
	assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode = coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_opcode;
	assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param = coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_param;
	assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size = coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_size;
	assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source = coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_source;
	assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink = coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_sink;
	assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied = coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_denied;
	assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data = coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_data;
	assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt = coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_corrupt;
	assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready = coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_ready;
	assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid = coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_valid;
	assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode = coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_opcode;
	assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param = coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_param;
	assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size = coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_size;
	assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink = coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_sink;
	assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied = coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_denied;
	assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data = coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_data;
	assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt = coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_corrupt;
	assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid = coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_valid;
	assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode = coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_opcode;
	assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param = coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_param;
	assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size = coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_size;
	assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source = coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_source;
	assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address = coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_address;
	assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask = coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_mask;
	assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data = coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_data;
	assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt = coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_corrupt;
	assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready = coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_ready;
	assign auto_fixedClockNode_out_1_clock = fixedClockNode_auto_out_2_clock;
	assign auto_fixedClockNode_out_1_reset = fixedClockNode_auto_out_2_reset;
	assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_clock = auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock;
	assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_reset = auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset;
	assign clockGroup_auto_in_member_subsystem_sbus_0_clock = subsystem_sbus_clock_groups_auto_out_member_subsystem_sbus_0_clock;
	assign clockGroup_auto_in_member_subsystem_sbus_0_reset = subsystem_sbus_clock_groups_auto_out_member_subsystem_sbus_0_reset;
	assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock;
	assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset;
	assign system_bus_xbar_clock = fixedClockNode_auto_out_0_clock;
	assign system_bus_xbar_reset = fixedClockNode_auto_out_0_reset;
	assign system_bus_xbar_auto_in_1_a_valid = fixer_auto_out_1_a_valid;
	assign system_bus_xbar_auto_in_1_a_bits_opcode = fixer_auto_out_1_a_bits_opcode;
	assign system_bus_xbar_auto_in_1_a_bits_param = fixer_auto_out_1_a_bits_param;
	assign system_bus_xbar_auto_in_1_a_bits_size = fixer_auto_out_1_a_bits_size;
	assign system_bus_xbar_auto_in_1_a_bits_source = fixer_auto_out_1_a_bits_source;
	assign system_bus_xbar_auto_in_1_a_bits_address = fixer_auto_out_1_a_bits_address;
	assign system_bus_xbar_auto_in_1_a_bits_mask = fixer_auto_out_1_a_bits_mask;
	assign system_bus_xbar_auto_in_1_a_bits_data = fixer_auto_out_1_a_bits_data;
	assign system_bus_xbar_auto_in_1_a_bits_corrupt = fixer_auto_out_1_a_bits_corrupt;
	assign system_bus_xbar_auto_in_1_d_ready = fixer_auto_out_1_d_ready;
	assign system_bus_xbar_auto_in_0_a_valid = fixer_auto_out_0_a_valid;
	assign system_bus_xbar_auto_in_0_a_bits_opcode = fixer_auto_out_0_a_bits_opcode;
	assign system_bus_xbar_auto_in_0_a_bits_param = fixer_auto_out_0_a_bits_param;
	assign system_bus_xbar_auto_in_0_a_bits_size = fixer_auto_out_0_a_bits_size;
	assign system_bus_xbar_auto_in_0_a_bits_source = fixer_auto_out_0_a_bits_source;
	assign system_bus_xbar_auto_in_0_a_bits_address = fixer_auto_out_0_a_bits_address;
	assign system_bus_xbar_auto_in_0_a_bits_mask = fixer_auto_out_0_a_bits_mask;
	assign system_bus_xbar_auto_in_0_a_bits_data = fixer_auto_out_0_a_bits_data;
	assign system_bus_xbar_auto_in_0_a_bits_corrupt = fixer_auto_out_0_a_bits_corrupt;
	assign system_bus_xbar_auto_in_0_d_ready = fixer_auto_out_0_d_ready;
	assign system_bus_xbar_auto_out_a_ready = coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_ready;
	assign system_bus_xbar_auto_out_d_valid = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_valid;
	assign system_bus_xbar_auto_out_d_bits_opcode = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_opcode;
	assign system_bus_xbar_auto_out_d_bits_param = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_param;
	assign system_bus_xbar_auto_out_d_bits_size = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_size;
	assign system_bus_xbar_auto_out_d_bits_source = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_source;
	assign system_bus_xbar_auto_out_d_bits_sink = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_sink;
	assign system_bus_xbar_auto_out_d_bits_denied = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_denied;
	assign system_bus_xbar_auto_out_d_bits_data = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_data;
	assign system_bus_xbar_auto_out_d_bits_corrupt = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_corrupt;
	assign fixer_clock = fixedClockNode_auto_out_0_clock;
	assign fixer_reset = fixedClockNode_auto_out_0_reset;
	assign fixer_auto_in_1_a_valid = coupler_from_tile_auto_tl_out_a_valid;
	assign fixer_auto_in_1_a_bits_opcode = coupler_from_tile_auto_tl_out_a_bits_opcode;
	assign fixer_auto_in_1_a_bits_param = coupler_from_tile_auto_tl_out_a_bits_param;
	assign fixer_auto_in_1_a_bits_size = coupler_from_tile_auto_tl_out_a_bits_size;
	assign fixer_auto_in_1_a_bits_source = coupler_from_tile_auto_tl_out_a_bits_source;
	assign fixer_auto_in_1_a_bits_address = coupler_from_tile_auto_tl_out_a_bits_address;
	assign fixer_auto_in_1_a_bits_mask = coupler_from_tile_auto_tl_out_a_bits_mask;
	assign fixer_auto_in_1_a_bits_data = coupler_from_tile_auto_tl_out_a_bits_data;
	assign fixer_auto_in_1_a_bits_corrupt = coupler_from_tile_auto_tl_out_a_bits_corrupt;
	assign fixer_auto_in_1_d_ready = coupler_from_tile_auto_tl_out_d_ready;
	assign fixer_auto_in_0_a_valid = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_valid;
	assign fixer_auto_in_0_a_bits_opcode = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_opcode;
	assign fixer_auto_in_0_a_bits_param = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_param;
	assign fixer_auto_in_0_a_bits_size = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_size;
	assign fixer_auto_in_0_a_bits_source = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_source;
	assign fixer_auto_in_0_a_bits_address = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_address;
	assign fixer_auto_in_0_a_bits_mask = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_mask;
	assign fixer_auto_in_0_a_bits_data = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_data;
	assign fixer_auto_in_0_a_bits_corrupt = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_corrupt;
	assign fixer_auto_in_0_d_ready = coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_ready;
	assign fixer_auto_out_1_a_ready = system_bus_xbar_auto_in_1_a_ready;
	assign fixer_auto_out_1_d_valid = system_bus_xbar_auto_in_1_d_valid;
	assign fixer_auto_out_1_d_bits_opcode = system_bus_xbar_auto_in_1_d_bits_opcode;
	assign fixer_auto_out_1_d_bits_param = system_bus_xbar_auto_in_1_d_bits_param;
	assign fixer_auto_out_1_d_bits_size = system_bus_xbar_auto_in_1_d_bits_size;
	assign fixer_auto_out_1_d_bits_source = system_bus_xbar_auto_in_1_d_bits_source;
	assign fixer_auto_out_1_d_bits_sink = system_bus_xbar_auto_in_1_d_bits_sink;
	assign fixer_auto_out_1_d_bits_denied = system_bus_xbar_auto_in_1_d_bits_denied;
	assign fixer_auto_out_1_d_bits_data = system_bus_xbar_auto_in_1_d_bits_data;
	assign fixer_auto_out_1_d_bits_corrupt = system_bus_xbar_auto_in_1_d_bits_corrupt;
	assign fixer_auto_out_0_a_ready = system_bus_xbar_auto_in_0_a_ready;
	assign fixer_auto_out_0_d_valid = system_bus_xbar_auto_in_0_d_valid;
	assign fixer_auto_out_0_d_bits_opcode = system_bus_xbar_auto_in_0_d_bits_opcode;
	assign fixer_auto_out_0_d_bits_param = system_bus_xbar_auto_in_0_d_bits_param;
	assign fixer_auto_out_0_d_bits_size = system_bus_xbar_auto_in_0_d_bits_size;
	assign fixer_auto_out_0_d_bits_sink = system_bus_xbar_auto_in_0_d_bits_sink;
	assign fixer_auto_out_0_d_bits_denied = system_bus_xbar_auto_in_0_d_bits_denied;
	assign fixer_auto_out_0_d_bits_data = system_bus_xbar_auto_in_0_d_bits_data;
	assign fixer_auto_out_0_d_bits_corrupt = system_bus_xbar_auto_in_0_d_bits_corrupt;
	assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_valid = system_bus_xbar_auto_out_a_valid;
	assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_opcode = system_bus_xbar_auto_out_a_bits_opcode;
	assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_param = system_bus_xbar_auto_out_a_bits_param;
	assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_size = system_bus_xbar_auto_out_a_bits_size;
	assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_source = system_bus_xbar_auto_out_a_bits_source;
	assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_address = system_bus_xbar_auto_out_a_bits_address;
	assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_mask = system_bus_xbar_auto_out_a_bits_mask;
	assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_data = system_bus_xbar_auto_out_a_bits_data;
	assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_corrupt = system_bus_xbar_auto_out_a_bits_corrupt;
	assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_ready = system_bus_xbar_auto_out_d_ready;
	assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_ready = auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready;
	assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_valid = auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid;
	assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_opcode = auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode;
	assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_param = auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param;
	assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_size = auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size;
	assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_source = auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source;
	assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_sink = auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink;
	assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_denied = auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied;
	assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_data = auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data;
	assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_corrupt = auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt;
	assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_ready = fixer_auto_in_0_a_ready;
	assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_valid = fixer_auto_in_0_d_valid;
	assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_opcode = fixer_auto_in_0_d_bits_opcode;
	assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_param = fixer_auto_in_0_d_bits_param;
	assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_size = fixer_auto_in_0_d_bits_size;
	assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_sink = fixer_auto_in_0_d_bits_sink;
	assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_denied = fixer_auto_in_0_d_bits_denied;
	assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_data = fixer_auto_in_0_d_bits_data;
	assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_corrupt = fixer_auto_in_0_d_bits_corrupt;
	assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_valid = auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid;
	assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_opcode = auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode;
	assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_param = auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param;
	assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_size = auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size;
	assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_source = auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source;
	assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_address = auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address;
	assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_mask = auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask;
	assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_data = auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data;
	assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_corrupt = auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_corrupt;
	assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_ready = auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready;
	assign coupler_from_tile_auto_tl_master_clock_xing_in_a_valid = auto_coupler_from_tile_tl_master_clock_xing_in_a_valid;
	assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_opcode = auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode;
	assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_param = auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param;
	assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_size = auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size;
	assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_source = auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source;
	assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_address = auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address;
	assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_mask = auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask;
	assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_data = auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data;
	assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_corrupt = auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_corrupt;
	assign coupler_from_tile_auto_tl_master_clock_xing_in_d_ready = auto_coupler_from_tile_tl_master_clock_xing_in_d_ready;
	assign coupler_from_tile_auto_tl_out_a_ready = fixer_auto_in_1_a_ready;
	assign coupler_from_tile_auto_tl_out_d_valid = fixer_auto_in_1_d_valid;
	assign coupler_from_tile_auto_tl_out_d_bits_opcode = fixer_auto_in_1_d_bits_opcode;
	assign coupler_from_tile_auto_tl_out_d_bits_param = fixer_auto_in_1_d_bits_param;
	assign coupler_from_tile_auto_tl_out_d_bits_size = fixer_auto_in_1_d_bits_size;
	assign coupler_from_tile_auto_tl_out_d_bits_source = fixer_auto_in_1_d_bits_source;
	assign coupler_from_tile_auto_tl_out_d_bits_sink = fixer_auto_in_1_d_bits_sink;
	assign coupler_from_tile_auto_tl_out_d_bits_denied = fixer_auto_in_1_d_bits_denied;
	assign coupler_from_tile_auto_tl_out_d_bits_data = fixer_auto_in_1_d_bits_data;
	assign coupler_from_tile_auto_tl_out_d_bits_corrupt = fixer_auto_in_1_d_bits_corrupt;
endmodule
module ClockGroupAggregator_1 (
	auto_in_member_subsystem_pbus_0_clock,
	auto_in_member_subsystem_pbus_0_reset,
	auto_out_member_subsystem_pbus_0_clock,
	auto_out_member_subsystem_pbus_0_reset
);
	input auto_in_member_subsystem_pbus_0_clock;
	input auto_in_member_subsystem_pbus_0_reset;
	output wire auto_out_member_subsystem_pbus_0_clock;
	output wire auto_out_member_subsystem_pbus_0_reset;
	assign auto_out_member_subsystem_pbus_0_clock = auto_in_member_subsystem_pbus_0_clock;
	assign auto_out_member_subsystem_pbus_0_reset = auto_in_member_subsystem_pbus_0_reset;
endmodule
module ClockGroup_1 (
	auto_in_member_subsystem_pbus_0_clock,
	auto_in_member_subsystem_pbus_0_reset,
	auto_out_clock,
	auto_out_reset
);
	input auto_in_member_subsystem_pbus_0_clock;
	input auto_in_member_subsystem_pbus_0_reset;
	output wire auto_out_clock;
	output wire auto_out_reset;
	assign auto_out_clock = auto_in_member_subsystem_pbus_0_clock;
	assign auto_out_reset = auto_in_member_subsystem_pbus_0_reset;
endmodule
module FixedClockBroadcast_1 (
	auto_in_clock,
	auto_in_reset,
	auto_out_1_clock,
	auto_out_1_reset,
	auto_out_0_clock,
	auto_out_0_reset
);
	input auto_in_clock;
	input auto_in_reset;
	output wire auto_out_1_clock;
	output wire auto_out_1_reset;
	output wire auto_out_0_clock;
	output wire auto_out_0_reset;
	assign auto_out_1_clock = auto_in_clock;
	assign auto_out_1_reset = auto_in_reset;
	assign auto_out_0_clock = auto_in_clock;
	assign auto_out_0_reset = auto_in_reset;
endmodule
module TLMonitor_4 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [30:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [30:0] _GEN_71 = {25'd0, is_aligned_mask};
	wire [30:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 31'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [30:0] _T_56 = io_in_a_bits_address ^ 31'h00004000;
	wire [31:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [31:0] _T_59 = $signed(_T_57) & -32'sh00001000;
	wire _T_60 = $signed(_T_59) == 32'sh00000000;
	wire [30:0] _T_61 = io_in_a_bits_address ^ 31'h00020000;
	wire [31:0] _T_62 = {1'b0, $signed(_T_61)};
	wire [31:0] _T_64 = $signed(_T_62) & -32'sh00010000;
	wire _T_65 = $signed(_T_64) == 32'sh00000000;
	wire [30:0] _T_66 = io_in_a_bits_address ^ 31'h10000000;
	wire [31:0] _T_67 = {1'b0, $signed(_T_66)};
	wire [31:0] _T_69 = $signed(_T_67) & -32'sh00001000;
	wire _T_70 = $signed(_T_69) == 32'sh00000000;
	wire [30:0] _T_71 = io_in_a_bits_address ^ 31'h54000000;
	wire [31:0] _T_72 = {1'b0, $signed(_T_71)};
	wire [31:0] _T_74 = $signed(_T_72) & -32'sh00001000;
	wire _T_75 = $signed(_T_74) == 32'sh00000000;
	wire _T_78 = ((_T_60 | _T_65) | _T_70) | _T_75;
	wire _T_128 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_132 = ~io_in_a_bits_mask;
	wire _T_133 = _T_132 == 4'h0;
	wire _T_137 = ~io_in_a_bits_corrupt;
	wire _T_141 = io_in_a_bits_opcode == 3'h7;
	wire _T_231 = io_in_a_bits_param != 3'h0;
	wire _T_244 = io_in_a_bits_opcode == 3'h4;
	wire _T_261 = io_in_a_bits_size <= 3'h6;
	wire _T_287 = _T_261 & _T_78;
	wire _T_298 = io_in_a_bits_param == 3'h0;
	wire _T_302 = io_in_a_bits_mask == mask;
	wire _T_310 = io_in_a_bits_opcode == 3'h0;
	wire _T_343 = (_T_60 | _T_70) | _T_75;
	wire _T_344 = _T_261 & _T_343;
	wire _T_354 = source_ok & _T_344;
	wire _T_372 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_430 = ~mask;
	wire [3:0] _T_431 = io_in_a_bits_mask & _T_430;
	wire _T_432 = _T_431 == 4'h0;
	wire _T_436 = io_in_a_bits_opcode == 3'h2;
	wire _T_485 = io_in_a_bits_param <= 3'h4;
	wire _T_493 = io_in_a_bits_opcode == 3'h3;
	wire _T_542 = io_in_a_bits_param <= 3'h3;
	wire _T_550 = io_in_a_bits_opcode == 3'h5;
	wire _T_599 = io_in_a_bits_param <= 3'h1;
	wire _T_611 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_615 = io_in_d_bits_opcode == 3'h6;
	wire _T_619 = io_in_d_bits_size >= 3'h2;
	wire _T_623 = io_in_d_bits_param == 2'h0;
	wire _T_627 = ~io_in_d_bits_corrupt;
	wire _T_631 = ~io_in_d_bits_denied;
	wire _T_635 = io_in_d_bits_opcode == 3'h4;
	wire _T_646 = io_in_d_bits_param <= 2'h2;
	wire _T_650 = io_in_d_bits_param != 2'h2;
	wire _T_663 = io_in_d_bits_opcode == 3'h5;
	wire _T_683 = _T_631 | io_in_d_bits_corrupt;
	wire _T_692 = io_in_d_bits_opcode == 3'h0;
	wire _T_709 = io_in_d_bits_opcode == 3'h1;
	wire _T_727 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [30:0] address;
	wire _T_757 = io_in_a_valid & ~a_first;
	wire _T_758 = io_in_a_bits_opcode == opcode;
	wire _T_762 = io_in_a_bits_param == param;
	wire _T_766 = io_in_a_bits_size == size;
	wire _T_770 = io_in_a_bits_source == source;
	wire _T_774 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_781 = io_in_d_valid & ~d_first;
	wire _T_782 = io_in_d_bits_opcode == opcode_1;
	wire _T_786 = io_in_d_bits_param == param_1;
	wire _T_790 = io_in_d_bits_size == size_1;
	wire _T_794 = io_in_d_bits_source == source_1;
	wire _T_798 = io_in_d_bits_sink == sink;
	wire _T_802 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_808 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire _T_811 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_813 = inflight >> io_in_a_bits_source;
	wire _T_815 = ~_T_813[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_819 = io_in_d_valid & d_first_1;
	wire _T_821 = ~_T_615;
	wire _T_822 = (io_in_d_valid & d_first_1) & ~_T_615;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_821 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_821 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_808 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_832 = inflight >> io_in_d_bits_source;
	wire _T_834 = _T_832[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_839 = io_in_d_bits_opcode == _GEN_40;
	wire _T_840 = (io_in_d_bits_opcode == _GEN_32) | _T_839;
	wire _T_844 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_851 = io_in_d_bits_opcode == _GEN_56;
	wire _T_852 = (io_in_d_bits_opcode == _GEN_48) | _T_851;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_856 = _GEN_82 == a_size_lookup;
	wire _T_866 = (((_T_819 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_821;
	wire _T_868 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_877 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_903 = (io_in_d_valid & d_first_2) & _T_615;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_615 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_615 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_911 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_921 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_941 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLFIFOFixer_1 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [30:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [30:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [30:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	TLMonitor_4 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_out_a_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid;
	assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_io_in_d_bits_param = auto_out_d_bits_param;
	assign monitor_io_in_d_bits_size = auto_out_d_bits_size;
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source;
	assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink;
	assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied;
	assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt;
endmodule
module TLXbar_1 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [30:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [30:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module TLMonitor_5 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [30:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [30:0] _GEN_71 = {25'd0, is_aligned_mask};
	wire [30:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 31'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [30:0] _T_56 = io_in_a_bits_address ^ 31'h00004000;
	wire [31:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [31:0] _T_59 = $signed(_T_57) & -32'sh00001000;
	wire _T_60 = $signed(_T_59) == 32'sh00000000;
	wire [30:0] _T_61 = io_in_a_bits_address ^ 31'h00020000;
	wire [31:0] _T_62 = {1'b0, $signed(_T_61)};
	wire [31:0] _T_64 = $signed(_T_62) & -32'sh00010000;
	wire _T_65 = $signed(_T_64) == 32'sh00000000;
	wire [30:0] _T_66 = io_in_a_bits_address ^ 31'h10000000;
	wire [31:0] _T_67 = {1'b0, $signed(_T_66)};
	wire [31:0] _T_69 = $signed(_T_67) & -32'sh00001000;
	wire _T_70 = $signed(_T_69) == 32'sh00000000;
	wire [30:0] _T_71 = io_in_a_bits_address ^ 31'h54000000;
	wire [31:0] _T_72 = {1'b0, $signed(_T_71)};
	wire [31:0] _T_74 = $signed(_T_72) & -32'sh00001000;
	wire _T_75 = $signed(_T_74) == 32'sh00000000;
	wire _T_78 = ((_T_60 | _T_65) | _T_70) | _T_75;
	wire _T_128 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_132 = ~io_in_a_bits_mask;
	wire _T_133 = _T_132 == 4'h0;
	wire _T_137 = ~io_in_a_bits_corrupt;
	wire _T_141 = io_in_a_bits_opcode == 3'h7;
	wire _T_231 = io_in_a_bits_param != 3'h0;
	wire _T_244 = io_in_a_bits_opcode == 3'h4;
	wire _T_261 = io_in_a_bits_size <= 3'h6;
	wire _T_287 = _T_261 & _T_78;
	wire _T_298 = io_in_a_bits_param == 3'h0;
	wire _T_302 = io_in_a_bits_mask == mask;
	wire _T_310 = io_in_a_bits_opcode == 3'h0;
	wire _T_343 = (_T_60 | _T_70) | _T_75;
	wire _T_344 = _T_261 & _T_343;
	wire _T_354 = source_ok & _T_344;
	wire _T_372 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_430 = ~mask;
	wire [3:0] _T_431 = io_in_a_bits_mask & _T_430;
	wire _T_432 = _T_431 == 4'h0;
	wire _T_436 = io_in_a_bits_opcode == 3'h2;
	wire _T_485 = io_in_a_bits_param <= 3'h4;
	wire _T_493 = io_in_a_bits_opcode == 3'h3;
	wire _T_542 = io_in_a_bits_param <= 3'h3;
	wire _T_550 = io_in_a_bits_opcode == 3'h5;
	wire _T_599 = io_in_a_bits_param <= 3'h1;
	wire _T_611 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_615 = io_in_d_bits_opcode == 3'h6;
	wire _T_619 = io_in_d_bits_size >= 3'h2;
	wire _T_623 = io_in_d_bits_param == 2'h0;
	wire _T_627 = ~io_in_d_bits_corrupt;
	wire _T_631 = ~io_in_d_bits_denied;
	wire _T_635 = io_in_d_bits_opcode == 3'h4;
	wire _T_646 = io_in_d_bits_param <= 2'h2;
	wire _T_650 = io_in_d_bits_param != 2'h2;
	wire _T_663 = io_in_d_bits_opcode == 3'h5;
	wire _T_683 = _T_631 | io_in_d_bits_corrupt;
	wire _T_692 = io_in_d_bits_opcode == 3'h0;
	wire _T_709 = io_in_d_bits_opcode == 3'h1;
	wire _T_727 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [30:0] address;
	wire _T_757 = io_in_a_valid & ~a_first;
	wire _T_758 = io_in_a_bits_opcode == opcode;
	wire _T_762 = io_in_a_bits_param == param;
	wire _T_766 = io_in_a_bits_size == size;
	wire _T_770 = io_in_a_bits_source == source;
	wire _T_774 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_781 = io_in_d_valid & ~d_first;
	wire _T_782 = io_in_d_bits_opcode == opcode_1;
	wire _T_786 = io_in_d_bits_param == param_1;
	wire _T_790 = io_in_d_bits_size == size_1;
	wire _T_794 = io_in_d_bits_source == source_1;
	wire _T_798 = io_in_d_bits_sink == sink;
	wire _T_802 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_808 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire _T_811 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_813 = inflight >> io_in_a_bits_source;
	wire _T_815 = ~_T_813[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_819 = io_in_d_valid & d_first_1;
	wire _T_821 = ~_T_615;
	wire _T_822 = (io_in_d_valid & d_first_1) & ~_T_615;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_821 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_821 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_808 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_832 = inflight >> io_in_d_bits_source;
	wire _T_834 = _T_832[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_839 = io_in_d_bits_opcode == _GEN_40;
	wire _T_840 = (io_in_d_bits_opcode == _GEN_32) | _T_839;
	wire _T_844 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_851 = io_in_d_bits_opcode == _GEN_56;
	wire _T_852 = (io_in_d_bits_opcode == _GEN_48) | _T_851;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_856 = _GEN_82 == a_size_lookup;
	wire _T_866 = (((_T_819 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_821;
	wire _T_868 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_877 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_903 = (io_in_d_valid & d_first_2) & _T_615;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_615 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_615 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_911 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_921 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_941 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLXbar_2 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_2_a_ready,
	auto_out_2_a_valid,
	auto_out_2_a_bits_opcode,
	auto_out_2_a_bits_param,
	auto_out_2_a_bits_size,
	auto_out_2_a_bits_source,
	auto_out_2_a_bits_address,
	auto_out_2_a_bits_mask,
	auto_out_2_a_bits_data,
	auto_out_2_a_bits_corrupt,
	auto_out_2_d_ready,
	auto_out_2_d_valid,
	auto_out_2_d_bits_opcode,
	auto_out_2_d_bits_size,
	auto_out_2_d_bits_source,
	auto_out_2_d_bits_data,
	auto_out_1_a_ready,
	auto_out_1_a_valid,
	auto_out_1_a_bits_opcode,
	auto_out_1_a_bits_param,
	auto_out_1_a_bits_size,
	auto_out_1_a_bits_source,
	auto_out_1_a_bits_address,
	auto_out_1_a_bits_mask,
	auto_out_1_a_bits_data,
	auto_out_1_a_bits_corrupt,
	auto_out_1_d_ready,
	auto_out_1_d_valid,
	auto_out_1_d_bits_opcode,
	auto_out_1_d_bits_param,
	auto_out_1_d_bits_size,
	auto_out_1_d_bits_source,
	auto_out_1_d_bits_sink,
	auto_out_1_d_bits_denied,
	auto_out_1_d_bits_data,
	auto_out_1_d_bits_corrupt,
	auto_out_0_a_ready,
	auto_out_0_a_valid,
	auto_out_0_a_bits_opcode,
	auto_out_0_a_bits_param,
	auto_out_0_a_bits_size,
	auto_out_0_a_bits_source,
	auto_out_0_a_bits_address,
	auto_out_0_a_bits_mask,
	auto_out_0_a_bits_data,
	auto_out_0_a_bits_corrupt,
	auto_out_0_d_ready,
	auto_out_0_d_valid,
	auto_out_0_d_bits_opcode,
	auto_out_0_d_bits_size,
	auto_out_0_d_bits_source,
	auto_out_0_d_bits_data
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [30:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_2_a_ready;
	output wire auto_out_2_a_valid;
	output wire [2:0] auto_out_2_a_bits_opcode;
	output wire [2:0] auto_out_2_a_bits_param;
	output wire [2:0] auto_out_2_a_bits_size;
	output wire [2:0] auto_out_2_a_bits_source;
	output wire [30:0] auto_out_2_a_bits_address;
	output wire [3:0] auto_out_2_a_bits_mask;
	output wire [31:0] auto_out_2_a_bits_data;
	output wire auto_out_2_a_bits_corrupt;
	output wire auto_out_2_d_ready;
	input auto_out_2_d_valid;
	input [2:0] auto_out_2_d_bits_opcode;
	input [2:0] auto_out_2_d_bits_size;
	input [2:0] auto_out_2_d_bits_source;
	input [31:0] auto_out_2_d_bits_data;
	input auto_out_1_a_ready;
	output wire auto_out_1_a_valid;
	output wire [2:0] auto_out_1_a_bits_opcode;
	output wire [2:0] auto_out_1_a_bits_param;
	output wire [2:0] auto_out_1_a_bits_size;
	output wire [2:0] auto_out_1_a_bits_source;
	output wire [28:0] auto_out_1_a_bits_address;
	output wire [3:0] auto_out_1_a_bits_mask;
	output wire [31:0] auto_out_1_a_bits_data;
	output wire auto_out_1_a_bits_corrupt;
	output wire auto_out_1_d_ready;
	input auto_out_1_d_valid;
	input [2:0] auto_out_1_d_bits_opcode;
	input [1:0] auto_out_1_d_bits_param;
	input [2:0] auto_out_1_d_bits_size;
	input [2:0] auto_out_1_d_bits_source;
	input auto_out_1_d_bits_sink;
	input auto_out_1_d_bits_denied;
	input [31:0] auto_out_1_d_bits_data;
	input auto_out_1_d_bits_corrupt;
	input auto_out_0_a_ready;
	output wire auto_out_0_a_valid;
	output wire [2:0] auto_out_0_a_bits_opcode;
	output wire [2:0] auto_out_0_a_bits_param;
	output wire [2:0] auto_out_0_a_bits_size;
	output wire [2:0] auto_out_0_a_bits_source;
	output wire [14:0] auto_out_0_a_bits_address;
	output wire [3:0] auto_out_0_a_bits_mask;
	output wire [31:0] auto_out_0_a_bits_data;
	output wire auto_out_0_a_bits_corrupt;
	output wire auto_out_0_d_ready;
	input auto_out_0_d_valid;
	input [2:0] auto_out_0_d_bits_opcode;
	input [2:0] auto_out_0_d_bits_size;
	input [2:0] auto_out_0_d_bits_source;
	input [31:0] auto_out_0_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [30:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	reg [3:0] beatsLeft;
	wire idle = beatsLeft == 4'h0;
	wire [2:0] readys_valid = {auto_out_2_d_valid, auto_out_1_d_valid, auto_out_0_d_valid};
	reg [2:0] readys_mask;
	wire [2:0] _readys_filter_T = ~readys_mask;
	wire [2:0] _readys_filter_T_1 = readys_valid & _readys_filter_T;
	wire [5:0] readys_filter = {_readys_filter_T_1, auto_out_2_d_valid, auto_out_1_d_valid, auto_out_0_d_valid};
	wire [5:0] _GEN_1 = {1'd0, readys_filter[5:1]};
	wire [5:0] _readys_unready_T_1 = readys_filter | _GEN_1;
	wire [5:0] _GEN_2 = {2'd0, _readys_unready_T_1[5:2]};
	wire [5:0] _readys_unready_T_3 = _readys_unready_T_1 | _GEN_2;
	wire [5:0] _readys_unready_T_6 = {readys_mask, 3'h0};
	wire [5:0] _GEN_3 = {1'd0, _readys_unready_T_3[5:1]};
	wire [5:0] readys_unready = _GEN_3 | _readys_unready_T_6;
	wire [2:0] _readys_readys_T_2 = readys_unready[5:3] & readys_unready[2:0];
	wire [2:0] readys_readys = ~_readys_readys_T_2;
	wire readys_0 = readys_readys[0];
	wire earlyWinner_0 = readys_0 & auto_out_0_d_valid;
	reg state_0;
	wire muxStateEarly_0 = (idle ? earlyWinner_0 : state_0);
	wire [2:0] _T_52 = (muxStateEarly_0 ? auto_out_0_d_bits_source : 3'h0);
	wire readys_1 = readys_readys[1];
	wire earlyWinner_1 = readys_1 & auto_out_1_d_valid;
	reg state_1;
	wire muxStateEarly_1 = (idle ? earlyWinner_1 : state_1);
	wire [2:0] _T_53 = (muxStateEarly_1 ? auto_out_1_d_bits_source : 3'h0);
	wire [2:0] _T_55 = _T_52 | _T_53;
	wire readys_2 = readys_readys[2];
	wire earlyWinner_2 = readys_2 & auto_out_2_d_valid;
	reg state_2;
	wire muxStateEarly_2 = (idle ? earlyWinner_2 : state_2);
	wire [2:0] _T_54 = (muxStateEarly_2 ? auto_out_2_d_bits_source : 3'h0);
	wire [31:0] _requestAIO_T_1 = {1'b0, $signed(auto_in_a_bits_address)};
	wire [31:0] _requestAIO_T_3 = $signed(_requestAIO_T_1) & 32'sh50020000;
	wire requestAIO_0_0 = $signed(_requestAIO_T_3) == 32'sh00000000;
	wire [30:0] _requestAIO_T_5 = auto_in_a_bits_address ^ 31'h00020000;
	wire [31:0] _requestAIO_T_6 = {1'b0, $signed(_requestAIO_T_5)};
	wire [31:0] _requestAIO_T_8 = $signed(_requestAIO_T_6) & 32'sh50020000;
	wire _requestAIO_T_9 = $signed(_requestAIO_T_8) == 32'sh00000000;
	wire [30:0] _requestAIO_T_10 = auto_in_a_bits_address ^ 31'h10000000;
	wire [31:0] _requestAIO_T_11 = {1'b0, $signed(_requestAIO_T_10)};
	wire [31:0] _requestAIO_T_13 = $signed(_requestAIO_T_11) & 32'sh50020000;
	wire _requestAIO_T_14 = $signed(_requestAIO_T_13) == 32'sh00000000;
	wire requestAIO_0_1 = _requestAIO_T_9 | _requestAIO_T_14;
	wire [30:0] _requestAIO_T_16 = auto_in_a_bits_address ^ 31'h50000000;
	wire [31:0] _requestAIO_T_17 = {1'b0, $signed(_requestAIO_T_16)};
	wire [31:0] _requestAIO_T_19 = $signed(_requestAIO_T_17) & 32'sh50020000;
	wire requestAIO_0_2 = $signed(_requestAIO_T_19) == 32'sh00000000;
	wire [12:0] _beatsDO_decode_T_1 = 13'h003f << auto_out_0_d_bits_size;
	wire [5:0] _beatsDO_decode_T_3 = ~_beatsDO_decode_T_1[5:0];
	wire [3:0] beatsDO_decode = _beatsDO_decode_T_3[5:2];
	wire beatsDO_opdata = auto_out_0_d_bits_opcode[0];
	wire [3:0] beatsDO_0 = (beatsDO_opdata ? beatsDO_decode : 4'h0);
	wire [12:0] _beatsDO_decode_T_5 = 13'h003f << auto_out_1_d_bits_size;
	wire [5:0] _beatsDO_decode_T_7 = ~_beatsDO_decode_T_5[5:0];
	wire [3:0] beatsDO_decode_1 = _beatsDO_decode_T_7[5:2];
	wire beatsDO_opdata_1 = auto_out_1_d_bits_opcode[0];
	wire [3:0] beatsDO_1 = (beatsDO_opdata_1 ? beatsDO_decode_1 : 4'h0);
	wire [12:0] _beatsDO_decode_T_9 = 13'h003f << auto_out_2_d_bits_size;
	wire [5:0] _beatsDO_decode_T_11 = ~_beatsDO_decode_T_9[5:0];
	wire [3:0] beatsDO_decode_2 = _beatsDO_decode_T_11[5:2];
	wire beatsDO_opdata_2 = auto_out_2_d_bits_opcode[0];
	wire [3:0] beatsDO_2 = (beatsDO_opdata_2 ? beatsDO_decode_2 : 4'h0);
	wire latch = idle & auto_in_d_ready;
	wire _readys_T_3 = ~reset;
	wire [2:0] _readys_mask_T = readys_readys & readys_valid;
	wire [3:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0};
	wire [2:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[2:0];
	wire [4:0] _readys_mask_T_4 = {_readys_mask_T_3, 2'h0};
	wire [2:0] _readys_mask_T_6 = _readys_mask_T_3 | _readys_mask_T_4[2:0];
	wire prefixOR_2 = earlyWinner_0 | earlyWinner_1;
	wire _prefixOR_T = prefixOR_2 | earlyWinner_2;
	wire _T_15 = (auto_out_0_d_valid | auto_out_1_d_valid) | auto_out_2_d_valid;
	wire _T_16 = ~((auto_out_0_d_valid | auto_out_1_d_valid) | auto_out_2_d_valid);
	wire [3:0] maskedBeats_0 = (earlyWinner_0 ? beatsDO_0 : 4'h0);
	wire [3:0] maskedBeats_1 = (earlyWinner_1 ? beatsDO_1 : 4'h0);
	wire [3:0] maskedBeats_2 = (earlyWinner_2 ? beatsDO_2 : 4'h0);
	wire [3:0] _initBeats_T = maskedBeats_0 | maskedBeats_1;
	wire [3:0] initBeats = _initBeats_T | maskedBeats_2;
	wire _sink_ACancel_earlyValid_T_6 = ((state_0 & auto_out_0_d_valid) | (state_1 & auto_out_1_d_valid)) | (state_2 & auto_out_2_d_valid);
	wire sink_ACancel_7_earlyValid = (idle ? _T_15 : _sink_ACancel_earlyValid_T_6);
	wire _beatsLeft_T_2 = auto_in_d_ready & sink_ACancel_7_earlyValid;
	wire [3:0] _GEN_4 = {3'd0, _beatsLeft_T_2};
	wire [3:0] _beatsLeft_T_4 = beatsLeft - _GEN_4;
	wire allowed_0 = (idle ? readys_0 : state_0);
	wire allowed_1 = (idle ? readys_1 : state_1);
	wire allowed_2 = (idle ? readys_2 : state_2);
	wire [31:0] _T_37 = (muxStateEarly_0 ? auto_out_0_d_bits_data : 32'h00000000);
	wire [31:0] _T_38 = (muxStateEarly_1 ? auto_out_1_d_bits_data : 32'h00000000);
	wire [31:0] _T_39 = (muxStateEarly_2 ? auto_out_2_d_bits_data : 32'h00000000);
	wire [31:0] _T_40 = _T_37 | _T_38;
	wire [2:0] _T_57 = (muxStateEarly_0 ? auto_out_0_d_bits_size : 3'h0);
	wire [2:0] _T_58 = (muxStateEarly_1 ? auto_out_1_d_bits_size : 3'h0);
	wire [2:0] _T_59 = (muxStateEarly_2 ? auto_out_2_d_bits_size : 3'h0);
	wire [2:0] _T_60 = _T_57 | _T_58;
	wire [2:0] _T_67 = (muxStateEarly_0 ? auto_out_0_d_bits_opcode : 3'h0);
	wire [2:0] _T_68 = (muxStateEarly_1 ? auto_out_1_d_bits_opcode : 3'h0);
	wire [2:0] _T_69 = (muxStateEarly_2 ? auto_out_2_d_bits_opcode : 3'h0);
	wire [2:0] _T_70 = _T_67 | _T_68;
	TLMonitor_5 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	assign auto_in_a_ready = ((requestAIO_0_0 & auto_out_0_a_ready) | (requestAIO_0_1 & auto_out_1_a_ready)) | (requestAIO_0_2 & auto_out_2_a_ready);
	assign auto_in_d_valid = (idle ? _T_15 : _sink_ACancel_earlyValid_T_6);
	assign auto_in_d_bits_opcode = _T_70 | _T_69;
	assign auto_in_d_bits_param = (muxStateEarly_1 ? auto_out_1_d_bits_param : 2'h0);
	assign auto_in_d_bits_size = _T_60 | _T_59;
	assign auto_in_d_bits_source = _T_55 | _T_54;
	assign auto_in_d_bits_sink = muxStateEarly_1 & auto_out_1_d_bits_sink;
	assign auto_in_d_bits_denied = muxStateEarly_1 & auto_out_1_d_bits_denied;
	assign auto_in_d_bits_data = _T_40 | _T_39;
	assign auto_in_d_bits_corrupt = muxStateEarly_1 & auto_out_1_d_bits_corrupt;
	assign auto_out_2_a_valid = auto_in_a_valid & requestAIO_0_2;
	assign auto_out_2_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_2_a_bits_param = auto_in_a_bits_param;
	assign auto_out_2_a_bits_size = auto_in_a_bits_size;
	assign auto_out_2_a_bits_source = auto_in_a_bits_source;
	assign auto_out_2_a_bits_address = auto_in_a_bits_address;
	assign auto_out_2_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_2_a_bits_data = auto_in_a_bits_data;
	assign auto_out_2_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_2_d_ready = auto_in_d_ready & allowed_2;
	assign auto_out_1_a_valid = auto_in_a_valid & requestAIO_0_1;
	assign auto_out_1_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_1_a_bits_param = auto_in_a_bits_param;
	assign auto_out_1_a_bits_size = auto_in_a_bits_size;
	assign auto_out_1_a_bits_source = auto_in_a_bits_source;
	assign auto_out_1_a_bits_address = auto_in_a_bits_address[28:0];
	assign auto_out_1_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_1_a_bits_data = auto_in_a_bits_data;
	assign auto_out_1_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_1_d_ready = auto_in_d_ready & allowed_1;
	assign auto_out_0_a_valid = auto_in_a_valid & requestAIO_0_0;
	assign auto_out_0_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_0_a_bits_param = auto_in_a_bits_param;
	assign auto_out_0_a_bits_size = auto_in_a_bits_size;
	assign auto_out_0_a_bits_source = auto_in_a_bits_source;
	assign auto_out_0_a_bits_address = auto_in_a_bits_address[14:0];
	assign auto_out_0_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_0_a_bits_data = auto_in_a_bits_data;
	assign auto_out_0_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_0_d_ready = auto_in_d_ready & allowed_0;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = ((requestAIO_0_0 & auto_out_0_a_ready) | (requestAIO_0_1 & auto_out_1_a_ready)) | (requestAIO_0_2 & auto_out_2_a_ready);
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = (idle ? _T_15 : _sink_ACancel_earlyValid_T_6);
	assign monitor_io_in_d_bits_opcode = _T_70 | _T_69;
	assign monitor_io_in_d_bits_param = (muxStateEarly_1 ? auto_out_1_d_bits_param : 2'h0);
	assign monitor_io_in_d_bits_size = _T_60 | _T_59;
	assign monitor_io_in_d_bits_source = _T_55 | _T_54;
	assign monitor_io_in_d_bits_sink = muxStateEarly_1 & auto_out_1_d_bits_sink;
	assign monitor_io_in_d_bits_denied = muxStateEarly_1 & auto_out_1_d_bits_denied;
	assign monitor_io_in_d_bits_corrupt = muxStateEarly_1 & auto_out_1_d_bits_corrupt;
	always @(posedge clock) begin
		if (reset)
			beatsLeft <= 4'h0;
		else if (latch)
			beatsLeft <= initBeats;
		else
			beatsLeft <= _beatsLeft_T_4;
		if (reset)
			readys_mask <= 3'h7;
		else if (latch & |readys_valid)
			readys_mask <= _readys_mask_T_6;
		if (reset)
			state_0 <= 1'h0;
		else if (idle)
			state_0 <= earlyWinner_0;
		if (reset)
			state_1 <= 1'h0;
		else if (idle)
			state_1 <= earlyWinner_1;
		if (reset)
			state_2 <= 1'h0;
		else if (idle)
			state_2 <= earlyWinner_2;
	end
endmodule
module TLMonitor_6 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [30:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [30:0] _GEN_71 = {25'd0, is_aligned_mask};
	wire [30:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 31'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [30:0] _T_56 = io_in_a_bits_address ^ 31'h00004000;
	wire [31:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [31:0] _T_59 = $signed(_T_57) & -32'sh00001000;
	wire _T_60 = $signed(_T_59) == 32'sh00000000;
	wire [30:0] _T_61 = io_in_a_bits_address ^ 31'h00020000;
	wire [31:0] _T_62 = {1'b0, $signed(_T_61)};
	wire [31:0] _T_64 = $signed(_T_62) & -32'sh00010000;
	wire _T_65 = $signed(_T_64) == 32'sh00000000;
	wire [30:0] _T_66 = io_in_a_bits_address ^ 31'h10000000;
	wire [31:0] _T_67 = {1'b0, $signed(_T_66)};
	wire [31:0] _T_69 = $signed(_T_67) & -32'sh00001000;
	wire _T_70 = $signed(_T_69) == 32'sh00000000;
	wire [30:0] _T_71 = io_in_a_bits_address ^ 31'h54000000;
	wire [31:0] _T_72 = {1'b0, $signed(_T_71)};
	wire [31:0] _T_74 = $signed(_T_72) & -32'sh00001000;
	wire _T_75 = $signed(_T_74) == 32'sh00000000;
	wire _T_78 = ((_T_60 | _T_65) | _T_70) | _T_75;
	wire _T_128 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_132 = ~io_in_a_bits_mask;
	wire _T_133 = _T_132 == 4'h0;
	wire _T_137 = ~io_in_a_bits_corrupt;
	wire _T_141 = io_in_a_bits_opcode == 3'h7;
	wire _T_231 = io_in_a_bits_param != 3'h0;
	wire _T_244 = io_in_a_bits_opcode == 3'h4;
	wire _T_261 = io_in_a_bits_size <= 3'h6;
	wire _T_287 = _T_261 & _T_78;
	wire _T_298 = io_in_a_bits_param == 3'h0;
	wire _T_302 = io_in_a_bits_mask == mask;
	wire _T_310 = io_in_a_bits_opcode == 3'h0;
	wire _T_343 = (_T_60 | _T_70) | _T_75;
	wire _T_344 = _T_261 & _T_343;
	wire _T_354 = source_ok & _T_344;
	wire _T_372 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_430 = ~mask;
	wire [3:0] _T_431 = io_in_a_bits_mask & _T_430;
	wire _T_432 = _T_431 == 4'h0;
	wire _T_436 = io_in_a_bits_opcode == 3'h2;
	wire _T_485 = io_in_a_bits_param <= 3'h4;
	wire _T_493 = io_in_a_bits_opcode == 3'h3;
	wire _T_542 = io_in_a_bits_param <= 3'h3;
	wire _T_550 = io_in_a_bits_opcode == 3'h5;
	wire _T_599 = io_in_a_bits_param <= 3'h1;
	wire _T_611 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_615 = io_in_d_bits_opcode == 3'h6;
	wire _T_619 = io_in_d_bits_size >= 3'h2;
	wire _T_623 = io_in_d_bits_param == 2'h0;
	wire _T_627 = ~io_in_d_bits_corrupt;
	wire _T_631 = ~io_in_d_bits_denied;
	wire _T_635 = io_in_d_bits_opcode == 3'h4;
	wire _T_646 = io_in_d_bits_param <= 2'h2;
	wire _T_650 = io_in_d_bits_param != 2'h2;
	wire _T_663 = io_in_d_bits_opcode == 3'h5;
	wire _T_683 = _T_631 | io_in_d_bits_corrupt;
	wire _T_692 = io_in_d_bits_opcode == 3'h0;
	wire _T_709 = io_in_d_bits_opcode == 3'h1;
	wire _T_727 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [30:0] address;
	wire _T_757 = io_in_a_valid & ~a_first;
	wire _T_758 = io_in_a_bits_opcode == opcode;
	wire _T_762 = io_in_a_bits_param == param;
	wire _T_766 = io_in_a_bits_size == size;
	wire _T_770 = io_in_a_bits_source == source;
	wire _T_774 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_781 = io_in_d_valid & ~d_first;
	wire _T_782 = io_in_d_bits_opcode == opcode_1;
	wire _T_786 = io_in_d_bits_param == param_1;
	wire _T_790 = io_in_d_bits_size == size_1;
	wire _T_794 = io_in_d_bits_source == source_1;
	wire _T_798 = io_in_d_bits_sink == sink;
	wire _T_802 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_808 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire [7:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire _T_811 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_813 = inflight >> io_in_a_bits_source;
	wire _T_815 = ~_T_813[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_819 = io_in_d_valid & d_first_1;
	wire _T_821 = ~_T_615;
	wire _T_822 = (io_in_d_valid & d_first_1) & ~_T_615;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [7:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_615 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_821 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_821 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_808 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_832 = inflight >> io_in_d_bits_source;
	wire _T_834 = _T_832[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_839 = io_in_d_bits_opcode == _GEN_40;
	wire _T_840 = (io_in_d_bits_opcode == _GEN_32) | _T_839;
	wire _T_844 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_851 = io_in_d_bits_opcode == _GEN_56;
	wire _T_852 = (io_in_d_bits_opcode == _GEN_48) | _T_851;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_856 = _GEN_82 == a_size_lookup;
	wire _T_866 = (((_T_819 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_821;
	wire _T_868 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set_wo_ready = _GEN_15[4:0];
	wire [4:0] d_clr_wo_ready = _GEN_21[4:0];
	wire _T_875 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_884 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_910 = (io_in_d_valid & d_first_2) & _T_615;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_615 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_615 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_918 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_928 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_953 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Queue (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_data,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [30:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input [31:0] io_enq_bits_data;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [30:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire [31:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg [2:0] ram_opcode [0:1];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [2:0] ram_param [0:1];
	wire ram_param_io_deq_bits_MPORT_en;
	wire ram_param_io_deq_bits_MPORT_addr;
	wire [2:0] ram_param_io_deq_bits_MPORT_data;
	wire [2:0] ram_param_MPORT_data;
	wire ram_param_MPORT_addr;
	wire ram_param_MPORT_mask;
	wire ram_param_MPORT_en;
	reg [2:0] ram_size [0:1];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [2:0] ram_size_io_deq_bits_MPORT_data;
	wire [2:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg [2:0] ram_source [0:1];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire [2:0] ram_source_io_deq_bits_MPORT_data;
	wire [2:0] ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg [30:0] ram_address [0:1];
	wire ram_address_io_deq_bits_MPORT_en;
	wire ram_address_io_deq_bits_MPORT_addr;
	wire [30:0] ram_address_io_deq_bits_MPORT_data;
	wire [30:0] ram_address_MPORT_data;
	wire ram_address_MPORT_addr;
	wire ram_address_MPORT_mask;
	wire ram_address_MPORT_en;
	reg [3:0] ram_mask [0:1];
	wire ram_mask_io_deq_bits_MPORT_en;
	wire ram_mask_io_deq_bits_MPORT_addr;
	wire [3:0] ram_mask_io_deq_bits_MPORT_data;
	wire [3:0] ram_mask_MPORT_data;
	wire ram_mask_MPORT_addr;
	wire ram_mask_MPORT_mask;
	wire ram_mask_MPORT_en;
	reg [31:0] ram_data [0:1];
	wire ram_data_io_deq_bits_MPORT_en;
	wire ram_data_io_deq_bits_MPORT_addr;
	wire [31:0] ram_data_io_deq_bits_MPORT_data;
	wire [31:0] ram_data_MPORT_data;
	wire ram_data_MPORT_addr;
	wire ram_data_MPORT_mask;
	wire ram_data_MPORT_en;
	reg ram_corrupt [0:1];
	wire ram_corrupt_io_deq_bits_MPORT_en;
	wire ram_corrupt_io_deq_bits_MPORT_addr;
	wire ram_corrupt_io_deq_bits_MPORT_data;
	wire ram_corrupt_MPORT_data;
	wire ram_corrupt_MPORT_addr;
	wire ram_corrupt_MPORT_mask;
	wire ram_corrupt_MPORT_en;
	reg value;
	reg value_1;
	reg maybe_full;
	wire ptr_match = value == value_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = value;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_param_io_deq_bits_MPORT_en = 1'h1;
	assign ram_param_io_deq_bits_MPORT_addr = value_1;
	assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr];
	assign ram_param_MPORT_data = io_enq_bits_param;
	assign ram_param_MPORT_addr = value;
	assign ram_param_MPORT_mask = 1'h1;
	assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = value_1;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = value;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = value_1;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = value;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_address_io_deq_bits_MPORT_en = 1'h1;
	assign ram_address_io_deq_bits_MPORT_addr = value_1;
	assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr];
	assign ram_address_MPORT_data = io_enq_bits_address;
	assign ram_address_MPORT_addr = value;
	assign ram_address_MPORT_mask = 1'h1;
	assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
	assign ram_mask_io_deq_bits_MPORT_addr = value_1;
	assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr];
	assign ram_mask_MPORT_data = io_enq_bits_mask;
	assign ram_mask_MPORT_addr = value;
	assign ram_mask_MPORT_mask = 1'h1;
	assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_data_io_deq_bits_MPORT_en = 1'h1;
	assign ram_data_io_deq_bits_MPORT_addr = value_1;
	assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr];
	assign ram_data_MPORT_data = io_enq_bits_data;
	assign ram_data_MPORT_addr = value;
	assign ram_data_MPORT_mask = 1'h1;
	assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
	assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
	assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr];
	assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
	assign ram_corrupt_MPORT_addr = value;
	assign ram_corrupt_MPORT_mask = 1'h1;
	assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data;
	assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data;
	assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data;
	assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_param_MPORT_en & ram_param_MPORT_mask)
			ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (ram_address_MPORT_en & ram_address_MPORT_mask)
			ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data;
		if (ram_mask_MPORT_en & ram_mask_MPORT_mask)
			ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data;
		if (ram_data_MPORT_en & ram_data_MPORT_mask)
			ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data;
		if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask)
			ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data;
		if (reset)
			value <= 1'h0;
		else if (do_enq)
			value <= value + 1'h1;
		if (reset)
			value_1 <= 1'h0;
		else if (do_deq)
			value_1 <= value_1 + 1'h1;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module Queue_1 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_sink,
	io_enq_bits_denied,
	io_enq_bits_data,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_sink,
	io_deq_bits_denied,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [1:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input io_enq_bits_sink;
	input io_enq_bits_denied;
	input [31:0] io_enq_bits_data;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [1:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire io_deq_bits_sink;
	output wire io_deq_bits_denied;
	output wire [31:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg [2:0] ram_opcode [0:1];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [1:0] ram_param [0:1];
	wire ram_param_io_deq_bits_MPORT_en;
	wire ram_param_io_deq_bits_MPORT_addr;
	wire [1:0] ram_param_io_deq_bits_MPORT_data;
	wire [1:0] ram_param_MPORT_data;
	wire ram_param_MPORT_addr;
	wire ram_param_MPORT_mask;
	wire ram_param_MPORT_en;
	reg [2:0] ram_size [0:1];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [2:0] ram_size_io_deq_bits_MPORT_data;
	wire [2:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg [2:0] ram_source [0:1];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire [2:0] ram_source_io_deq_bits_MPORT_data;
	wire [2:0] ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg ram_sink [0:1];
	wire ram_sink_io_deq_bits_MPORT_en;
	wire ram_sink_io_deq_bits_MPORT_addr;
	wire ram_sink_io_deq_bits_MPORT_data;
	wire ram_sink_MPORT_data;
	wire ram_sink_MPORT_addr;
	wire ram_sink_MPORT_mask;
	wire ram_sink_MPORT_en;
	reg ram_denied [0:1];
	wire ram_denied_io_deq_bits_MPORT_en;
	wire ram_denied_io_deq_bits_MPORT_addr;
	wire ram_denied_io_deq_bits_MPORT_data;
	wire ram_denied_MPORT_data;
	wire ram_denied_MPORT_addr;
	wire ram_denied_MPORT_mask;
	wire ram_denied_MPORT_en;
	reg [31:0] ram_data [0:1];
	wire ram_data_io_deq_bits_MPORT_en;
	wire ram_data_io_deq_bits_MPORT_addr;
	wire [31:0] ram_data_io_deq_bits_MPORT_data;
	wire [31:0] ram_data_MPORT_data;
	wire ram_data_MPORT_addr;
	wire ram_data_MPORT_mask;
	wire ram_data_MPORT_en;
	reg ram_corrupt [0:1];
	wire ram_corrupt_io_deq_bits_MPORT_en;
	wire ram_corrupt_io_deq_bits_MPORT_addr;
	wire ram_corrupt_io_deq_bits_MPORT_data;
	wire ram_corrupt_MPORT_data;
	wire ram_corrupt_MPORT_addr;
	wire ram_corrupt_MPORT_mask;
	wire ram_corrupt_MPORT_en;
	reg value;
	reg value_1;
	reg maybe_full;
	wire ptr_match = value == value_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = value;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_param_io_deq_bits_MPORT_en = 1'h1;
	assign ram_param_io_deq_bits_MPORT_addr = value_1;
	assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr];
	assign ram_param_MPORT_data = io_enq_bits_param;
	assign ram_param_MPORT_addr = value;
	assign ram_param_MPORT_mask = 1'h1;
	assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = value_1;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = value;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = value_1;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = value;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_sink_io_deq_bits_MPORT_en = 1'h1;
	assign ram_sink_io_deq_bits_MPORT_addr = value_1;
	assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr];
	assign ram_sink_MPORT_data = io_enq_bits_sink;
	assign ram_sink_MPORT_addr = value;
	assign ram_sink_MPORT_mask = 1'h1;
	assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_denied_io_deq_bits_MPORT_en = 1'h1;
	assign ram_denied_io_deq_bits_MPORT_addr = value_1;
	assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr];
	assign ram_denied_MPORT_data = io_enq_bits_denied;
	assign ram_denied_MPORT_addr = value;
	assign ram_denied_MPORT_mask = 1'h1;
	assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_data_io_deq_bits_MPORT_en = 1'h1;
	assign ram_data_io_deq_bits_MPORT_addr = value_1;
	assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr];
	assign ram_data_MPORT_data = io_enq_bits_data;
	assign ram_data_MPORT_addr = value;
	assign ram_data_MPORT_mask = 1'h1;
	assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
	assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
	assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr];
	assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
	assign ram_corrupt_MPORT_addr = value;
	assign ram_corrupt_MPORT_mask = 1'h1;
	assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data;
	assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data;
	assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data;
	assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_param_MPORT_en & ram_param_MPORT_mask)
			ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (ram_sink_MPORT_en & ram_sink_MPORT_mask)
			ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data;
		if (ram_denied_MPORT_en & ram_denied_MPORT_mask)
			ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data;
		if (ram_data_MPORT_en & ram_data_MPORT_mask)
			ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data;
		if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask)
			ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data;
		if (reset)
			value <= 1'h0;
		else if (do_enq)
			value <= value + 1'h1;
		if (reset)
			value_1 <= 1'h0;
		else if (do_deq)
			value_1 <= value_1 + 1'h1;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module TLBuffer_1 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [30:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [30:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [30:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire bundleOut_0_a_q_clock;
	wire bundleOut_0_a_q_reset;
	wire bundleOut_0_a_q_io_enq_ready;
	wire bundleOut_0_a_q_io_enq_valid;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_param;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_size;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_source;
	wire [30:0] bundleOut_0_a_q_io_enq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_data;
	wire bundleOut_0_a_q_io_enq_bits_corrupt;
	wire bundleOut_0_a_q_io_deq_ready;
	wire bundleOut_0_a_q_io_deq_valid;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_param;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_size;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_source;
	wire [30:0] bundleOut_0_a_q_io_deq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_data;
	wire bundleOut_0_a_q_io_deq_bits_corrupt;
	wire bundleIn_0_d_q_clock;
	wire bundleIn_0_d_q_reset;
	wire bundleIn_0_d_q_io_enq_ready;
	wire bundleIn_0_d_q_io_enq_valid;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_enq_bits_param;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_size;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_source;
	wire bundleIn_0_d_q_io_enq_bits_sink;
	wire bundleIn_0_d_q_io_enq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_enq_bits_data;
	wire bundleIn_0_d_q_io_enq_bits_corrupt;
	wire bundleIn_0_d_q_io_deq_ready;
	wire bundleIn_0_d_q_io_deq_valid;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_param;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_size;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_source;
	wire bundleIn_0_d_q_io_deq_bits_sink;
	wire bundleIn_0_d_q_io_deq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_deq_bits_data;
	wire bundleIn_0_d_q_io_deq_bits_corrupt;
	TLMonitor_6 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Queue bundleOut_0_a_q(
		.clock(bundleOut_0_a_q_clock),
		.reset(bundleOut_0_a_q_reset),
		.io_enq_ready(bundleOut_0_a_q_io_enq_ready),
		.io_enq_valid(bundleOut_0_a_q_io_enq_valid),
		.io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
		.io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
		.io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
		.io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
		.io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
		.io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleOut_0_a_q_io_deq_ready),
		.io_deq_valid(bundleOut_0_a_q_io_deq_valid),
		.io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
		.io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
		.io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
		.io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
		.io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
		.io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
	);
	Queue_1 bundleIn_0_d_q(
		.clock(bundleIn_0_d_q_clock),
		.reset(bundleIn_0_d_q_reset),
		.io_enq_ready(bundleIn_0_d_q_io_enq_ready),
		.io_enq_valid(bundleIn_0_d_q_io_enq_valid),
		.io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
		.io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
		.io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
		.io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
		.io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
		.io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleIn_0_d_q_io_deq_ready),
		.io_deq_valid(bundleIn_0_d_q_io_deq_valid),
		.io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
		.io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
		.io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
		.io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
		.io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
		.io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data;
	assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid;
	assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode;
	assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param;
	assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size;
	assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source;
	assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address;
	assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask;
	assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data;
	assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt;
	assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign bundleOut_0_a_q_clock = clock;
	assign bundleOut_0_a_q_reset = reset;
	assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid;
	assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param;
	assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size;
	assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source;
	assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address;
	assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask;
	assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data;
	assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready;
	assign bundleIn_0_d_q_clock = clock;
	assign bundleIn_0_d_q_reset = reset;
	assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid;
	assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign bundleIn_0_d_q_io_enq_bits_param = auto_out_d_bits_param;
	assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size;
	assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source;
	assign bundleIn_0_d_q_io_enq_bits_sink = auto_out_d_bits_sink;
	assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied;
	assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data;
	assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt;
	assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready;
endmodule
module TLMonitor_7 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [30:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [30:0] _GEN_71 = {25'd0, is_aligned_mask};
	wire [30:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 31'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [30:0] _T_56 = io_in_a_bits_address ^ 31'h00004000;
	wire [31:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [31:0] _T_59 = $signed(_T_57) & -32'sh00001000;
	wire _T_60 = $signed(_T_59) == 32'sh00000000;
	wire [30:0] _T_61 = io_in_a_bits_address ^ 31'h00020000;
	wire [31:0] _T_62 = {1'b0, $signed(_T_61)};
	wire [31:0] _T_64 = $signed(_T_62) & -32'sh00010000;
	wire _T_65 = $signed(_T_64) == 32'sh00000000;
	wire [30:0] _T_66 = io_in_a_bits_address ^ 31'h10000000;
	wire [31:0] _T_67 = {1'b0, $signed(_T_66)};
	wire [31:0] _T_69 = $signed(_T_67) & -32'sh00001000;
	wire _T_70 = $signed(_T_69) == 32'sh00000000;
	wire [30:0] _T_71 = io_in_a_bits_address ^ 31'h54000000;
	wire [31:0] _T_72 = {1'b0, $signed(_T_71)};
	wire [31:0] _T_74 = $signed(_T_72) & -32'sh00001000;
	wire _T_75 = $signed(_T_74) == 32'sh00000000;
	wire _T_78 = ((_T_60 | _T_65) | _T_70) | _T_75;
	wire _T_128 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_132 = ~io_in_a_bits_mask;
	wire _T_133 = _T_132 == 4'h0;
	wire _T_137 = ~io_in_a_bits_corrupt;
	wire _T_141 = io_in_a_bits_opcode == 3'h7;
	wire _T_231 = io_in_a_bits_param != 3'h0;
	wire _T_244 = io_in_a_bits_opcode == 3'h4;
	wire _T_261 = io_in_a_bits_size <= 3'h6;
	wire _T_287 = _T_261 & _T_78;
	wire _T_298 = io_in_a_bits_param == 3'h0;
	wire _T_302 = io_in_a_bits_mask == mask;
	wire _T_310 = io_in_a_bits_opcode == 3'h0;
	wire _T_343 = (_T_60 | _T_70) | _T_75;
	wire _T_344 = _T_261 & _T_343;
	wire _T_354 = source_ok & _T_344;
	wire _T_372 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_430 = ~mask;
	wire [3:0] _T_431 = io_in_a_bits_mask & _T_430;
	wire _T_432 = _T_431 == 4'h0;
	wire _T_436 = io_in_a_bits_opcode == 3'h2;
	wire _T_450 = io_in_a_bits_size <= 3'h2;
	wire _T_470 = _T_450 & _T_343;
	wire _T_480 = source_ok & _T_470;
	wire _T_490 = io_in_a_bits_param <= 3'h4;
	wire _T_498 = io_in_a_bits_opcode == 3'h3;
	wire _T_552 = io_in_a_bits_param <= 3'h3;
	wire _T_560 = io_in_a_bits_opcode == 3'h5;
	wire _T_609 = io_in_a_bits_param <= 3'h1;
	wire _T_621 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_625 = io_in_d_bits_opcode == 3'h6;
	wire _T_629 = io_in_d_bits_size >= 3'h2;
	wire _T_633 = io_in_d_bits_param == 2'h0;
	wire _T_637 = ~io_in_d_bits_corrupt;
	wire _T_641 = ~io_in_d_bits_denied;
	wire _T_645 = io_in_d_bits_opcode == 3'h4;
	wire _T_656 = io_in_d_bits_param <= 2'h2;
	wire _T_660 = io_in_d_bits_param != 2'h2;
	wire _T_673 = io_in_d_bits_opcode == 3'h5;
	wire _T_693 = _T_641 | io_in_d_bits_corrupt;
	wire _T_702 = io_in_d_bits_opcode == 3'h0;
	wire _T_719 = io_in_d_bits_opcode == 3'h1;
	wire _T_737 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [30:0] address;
	wire _T_767 = io_in_a_valid & ~a_first;
	wire _T_768 = io_in_a_bits_opcode == opcode;
	wire _T_772 = io_in_a_bits_param == param;
	wire _T_776 = io_in_a_bits_size == size;
	wire _T_780 = io_in_a_bits_source == source;
	wire _T_784 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_791 = io_in_d_valid & ~d_first;
	wire _T_792 = io_in_d_bits_opcode == opcode_1;
	wire _T_796 = io_in_d_bits_param == param_1;
	wire _T_800 = io_in_d_bits_size == size_1;
	wire _T_804 = io_in_d_bits_source == source_1;
	wire _T_808 = io_in_d_bits_sink == sink;
	wire _T_812 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_818 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire [7:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire _T_821 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_823 = inflight >> io_in_a_bits_source;
	wire _T_825 = ~_T_823[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_829 = io_in_d_valid & d_first_1;
	wire _T_831 = ~_T_625;
	wire _T_832 = (io_in_d_valid & d_first_1) & ~_T_625;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [7:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_625 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_831 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_831 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_818 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_842 = inflight >> io_in_d_bits_source;
	wire _T_844 = _T_842[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_849 = io_in_d_bits_opcode == _GEN_40;
	wire _T_850 = (io_in_d_bits_opcode == _GEN_32) | _T_849;
	wire _T_854 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_861 = io_in_d_bits_opcode == _GEN_56;
	wire _T_862 = (io_in_d_bits_opcode == _GEN_48) | _T_861;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_866 = _GEN_82 == a_size_lookup;
	wire _T_876 = (((_T_829 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_831;
	wire _T_878 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set_wo_ready = _GEN_15[4:0];
	wire [4:0] d_clr_wo_ready = _GEN_21[4:0];
	wire _T_885 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_894 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_920 = (io_in_d_valid & d_first_2) & _T_625;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_625 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_625 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_928 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_938 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_963 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLAtomicAutomata (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [30:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [30:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [30:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	reg [1:0] cam_s_0_state;
	reg [2:0] cam_a_0_bits_opcode;
	reg [2:0] cam_a_0_bits_param;
	reg [2:0] cam_a_0_bits_size;
	reg [2:0] cam_a_0_bits_source;
	reg [30:0] cam_a_0_bits_address;
	reg [3:0] cam_a_0_bits_mask;
	reg [31:0] cam_a_0_bits_data;
	reg cam_a_0_bits_corrupt;
	reg [3:0] cam_a_0_lut;
	reg [31:0] cam_d_0_data;
	reg cam_d_0_denied;
	reg cam_d_0_corrupt;
	wire cam_free_0 = cam_s_0_state == 2'h0;
	wire cam_amo_0 = cam_s_0_state == 2'h2;
	wire cam_abusy_0 = (cam_s_0_state == 2'h3) | cam_amo_0;
	wire cam_dmatch_0 = cam_s_0_state != 2'h0;
	wire a_isLogical = auto_in_a_bits_opcode == 3'h3;
	wire a_isArithmetic = auto_in_a_bits_opcode == 3'h2;
	wire _a_isSupported_T = (a_isArithmetic ? 1'h0 : 1'h1);
	wire a_isSupported = (a_isLogical ? 1'h0 : _a_isSupported_T);
	wire [1:0] indexes_0 = {cam_a_0_bits_data[0], cam_d_0_data[0]};
	wire [1:0] indexes_1 = {cam_a_0_bits_data[1], cam_d_0_data[1]};
	wire [1:0] indexes_2 = {cam_a_0_bits_data[2], cam_d_0_data[2]};
	wire [1:0] indexes_3 = {cam_a_0_bits_data[3], cam_d_0_data[3]};
	wire [1:0] indexes_4 = {cam_a_0_bits_data[4], cam_d_0_data[4]};
	wire [1:0] indexes_5 = {cam_a_0_bits_data[5], cam_d_0_data[5]};
	wire [1:0] indexes_6 = {cam_a_0_bits_data[6], cam_d_0_data[6]};
	wire [1:0] indexes_7 = {cam_a_0_bits_data[7], cam_d_0_data[7]};
	wire [1:0] indexes_8 = {cam_a_0_bits_data[8], cam_d_0_data[8]};
	wire [1:0] indexes_9 = {cam_a_0_bits_data[9], cam_d_0_data[9]};
	wire [1:0] indexes_10 = {cam_a_0_bits_data[10], cam_d_0_data[10]};
	wire [1:0] indexes_11 = {cam_a_0_bits_data[11], cam_d_0_data[11]};
	wire [1:0] indexes_12 = {cam_a_0_bits_data[12], cam_d_0_data[12]};
	wire [1:0] indexes_13 = {cam_a_0_bits_data[13], cam_d_0_data[13]};
	wire [1:0] indexes_14 = {cam_a_0_bits_data[14], cam_d_0_data[14]};
	wire [1:0] indexes_15 = {cam_a_0_bits_data[15], cam_d_0_data[15]};
	wire [1:0] indexes_16 = {cam_a_0_bits_data[16], cam_d_0_data[16]};
	wire [1:0] indexes_17 = {cam_a_0_bits_data[17], cam_d_0_data[17]};
	wire [1:0] indexes_18 = {cam_a_0_bits_data[18], cam_d_0_data[18]};
	wire [1:0] indexes_19 = {cam_a_0_bits_data[19], cam_d_0_data[19]};
	wire [1:0] indexes_20 = {cam_a_0_bits_data[20], cam_d_0_data[20]};
	wire [1:0] indexes_21 = {cam_a_0_bits_data[21], cam_d_0_data[21]};
	wire [1:0] indexes_22 = {cam_a_0_bits_data[22], cam_d_0_data[22]};
	wire [1:0] indexes_23 = {cam_a_0_bits_data[23], cam_d_0_data[23]};
	wire [1:0] indexes_24 = {cam_a_0_bits_data[24], cam_d_0_data[24]};
	wire [1:0] indexes_25 = {cam_a_0_bits_data[25], cam_d_0_data[25]};
	wire [1:0] indexes_26 = {cam_a_0_bits_data[26], cam_d_0_data[26]};
	wire [1:0] indexes_27 = {cam_a_0_bits_data[27], cam_d_0_data[27]};
	wire [1:0] indexes_28 = {cam_a_0_bits_data[28], cam_d_0_data[28]};
	wire [1:0] indexes_29 = {cam_a_0_bits_data[29], cam_d_0_data[29]};
	wire [1:0] indexes_30 = {cam_a_0_bits_data[30], cam_d_0_data[30]};
	wire [1:0] indexes_31 = {cam_a_0_bits_data[31], cam_d_0_data[31]};
	wire [3:0] _logic_out_T = cam_a_0_lut >> indexes_0;
	wire [3:0] _logic_out_T_2 = cam_a_0_lut >> indexes_1;
	wire [3:0] _logic_out_T_4 = cam_a_0_lut >> indexes_2;
	wire [3:0] _logic_out_T_6 = cam_a_0_lut >> indexes_3;
	wire [3:0] _logic_out_T_8 = cam_a_0_lut >> indexes_4;
	wire [3:0] _logic_out_T_10 = cam_a_0_lut >> indexes_5;
	wire [3:0] _logic_out_T_12 = cam_a_0_lut >> indexes_6;
	wire [3:0] _logic_out_T_14 = cam_a_0_lut >> indexes_7;
	wire [3:0] _logic_out_T_16 = cam_a_0_lut >> indexes_8;
	wire [3:0] _logic_out_T_18 = cam_a_0_lut >> indexes_9;
	wire [3:0] _logic_out_T_20 = cam_a_0_lut >> indexes_10;
	wire [3:0] _logic_out_T_22 = cam_a_0_lut >> indexes_11;
	wire [3:0] _logic_out_T_24 = cam_a_0_lut >> indexes_12;
	wire [3:0] _logic_out_T_26 = cam_a_0_lut >> indexes_13;
	wire [3:0] _logic_out_T_28 = cam_a_0_lut >> indexes_14;
	wire [3:0] _logic_out_T_30 = cam_a_0_lut >> indexes_15;
	wire [3:0] _logic_out_T_32 = cam_a_0_lut >> indexes_16;
	wire [3:0] _logic_out_T_34 = cam_a_0_lut >> indexes_17;
	wire [3:0] _logic_out_T_36 = cam_a_0_lut >> indexes_18;
	wire [3:0] _logic_out_T_38 = cam_a_0_lut >> indexes_19;
	wire [3:0] _logic_out_T_40 = cam_a_0_lut >> indexes_20;
	wire [3:0] _logic_out_T_42 = cam_a_0_lut >> indexes_21;
	wire [3:0] _logic_out_T_44 = cam_a_0_lut >> indexes_22;
	wire [3:0] _logic_out_T_46 = cam_a_0_lut >> indexes_23;
	wire [3:0] _logic_out_T_48 = cam_a_0_lut >> indexes_24;
	wire [3:0] _logic_out_T_50 = cam_a_0_lut >> indexes_25;
	wire [3:0] _logic_out_T_52 = cam_a_0_lut >> indexes_26;
	wire [3:0] _logic_out_T_54 = cam_a_0_lut >> indexes_27;
	wire [3:0] _logic_out_T_56 = cam_a_0_lut >> indexes_28;
	wire [3:0] _logic_out_T_58 = cam_a_0_lut >> indexes_29;
	wire [3:0] _logic_out_T_60 = cam_a_0_lut >> indexes_30;
	wire [3:0] _logic_out_T_62 = cam_a_0_lut >> indexes_31;
	wire [7:0] logic_out_lo_lo = {_logic_out_T_14[0], _logic_out_T_12[0], _logic_out_T_10[0], _logic_out_T_8[0], _logic_out_T_6[0], _logic_out_T_4[0], _logic_out_T_2[0], _logic_out_T[0]};
	wire [15:0] logic_out_lo = {_logic_out_T_30[0], _logic_out_T_28[0], _logic_out_T_26[0], _logic_out_T_24[0], _logic_out_T_22[0], _logic_out_T_20[0], _logic_out_T_18[0], _logic_out_T_16[0], logic_out_lo_lo};
	wire [7:0] logic_out_hi_lo = {_logic_out_T_46[0], _logic_out_T_44[0], _logic_out_T_42[0], _logic_out_T_40[0], _logic_out_T_38[0], _logic_out_T_36[0], _logic_out_T_34[0], _logic_out_T_32[0]};
	wire [31:0] logic_out = {_logic_out_T_62[0], _logic_out_T_60[0], _logic_out_T_58[0], _logic_out_T_56[0], _logic_out_T_54[0], _logic_out_T_52[0], _logic_out_T_50[0], _logic_out_T_48[0], logic_out_hi_lo, logic_out_lo};
	wire unsigned_ = cam_a_0_bits_param[1];
	wire take_max = cam_a_0_bits_param[0];
	wire adder = cam_a_0_bits_param[2];
	wire [3:0] _signSel_T = ~cam_a_0_bits_mask;
	wire [3:0] _GEN_39 = {1'd0, cam_a_0_bits_mask[3:1]};
	wire [3:0] _signSel_T_2 = _signSel_T | _GEN_39;
	wire [3:0] signSel = ~_signSel_T_2;
	wire [3:0] signbits_a = {cam_a_0_bits_data[31], cam_a_0_bits_data[23], cam_a_0_bits_data[15], cam_a_0_bits_data[7]};
	wire [3:0] signbits_d = {cam_d_0_data[31], cam_d_0_data[23], cam_d_0_data[15], cam_d_0_data[7]};
	wire [3:0] _signbit_a_T = signbits_a & signSel;
	wire [4:0] _signbit_a_T_1 = {_signbit_a_T, 1'h0};
	wire [3:0] signbit_a = _signbit_a_T_1[3:0];
	wire [3:0] _signbit_d_T = signbits_d & signSel;
	wire [4:0] _signbit_d_T_1 = {_signbit_d_T, 1'h0};
	wire [3:0] signbit_d = _signbit_d_T_1[3:0];
	wire [4:0] _signext_a_T = {signbit_a, 1'h0};
	wire [3:0] _signext_a_T_2 = signbit_a | _signext_a_T[3:0];
	wire [5:0] _signext_a_T_3 = {_signext_a_T_2, 2'h0};
	wire [3:0] _signext_a_T_5 = _signext_a_T_2 | _signext_a_T_3[3:0];
	wire [7:0] _signext_a_T_12 = (_signext_a_T_5[0] ? 8'hff : 8'h00);
	wire [7:0] _signext_a_T_14 = (_signext_a_T_5[1] ? 8'hff : 8'h00);
	wire [7:0] _signext_a_T_16 = (_signext_a_T_5[2] ? 8'hff : 8'h00);
	wire [7:0] _signext_a_T_18 = (_signext_a_T_5[3] ? 8'hff : 8'h00);
	wire [31:0] signext_a = {_signext_a_T_18, _signext_a_T_16, _signext_a_T_14, _signext_a_T_12};
	wire [4:0] _signext_d_T = {signbit_d, 1'h0};
	wire [3:0] _signext_d_T_2 = signbit_d | _signext_d_T[3:0];
	wire [5:0] _signext_d_T_3 = {_signext_d_T_2, 2'h0};
	wire [3:0] _signext_d_T_5 = _signext_d_T_2 | _signext_d_T_3[3:0];
	wire [7:0] _signext_d_T_12 = (_signext_d_T_5[0] ? 8'hff : 8'h00);
	wire [7:0] _signext_d_T_14 = (_signext_d_T_5[1] ? 8'hff : 8'h00);
	wire [7:0] _signext_d_T_16 = (_signext_d_T_5[2] ? 8'hff : 8'h00);
	wire [7:0] _signext_d_T_18 = (_signext_d_T_5[3] ? 8'hff : 8'h00);
	wire [31:0] signext_d = {_signext_d_T_18, _signext_d_T_16, _signext_d_T_14, _signext_d_T_12};
	wire [7:0] _wide_mask_T_5 = (cam_a_0_bits_mask[0] ? 8'hff : 8'h00);
	wire [7:0] _wide_mask_T_7 = (cam_a_0_bits_mask[1] ? 8'hff : 8'h00);
	wire [7:0] _wide_mask_T_9 = (cam_a_0_bits_mask[2] ? 8'hff : 8'h00);
	wire [7:0] _wide_mask_T_11 = (cam_a_0_bits_mask[3] ? 8'hff : 8'h00);
	wire [31:0] wide_mask = {_wide_mask_T_11, _wide_mask_T_9, _wide_mask_T_7, _wide_mask_T_5};
	wire [31:0] _a_a_ext_T = cam_a_0_bits_data & wide_mask;
	wire [31:0] a_a_ext = _a_a_ext_T | signext_a;
	wire [31:0] _a_d_ext_T = cam_d_0_data & wide_mask;
	wire [31:0] a_d_ext = _a_d_ext_T | signext_d;
	wire [31:0] _a_d_inv_T = ~a_d_ext;
	wire [31:0] a_d_inv = (adder ? a_d_ext : _a_d_inv_T);
	wire [31:0] adder_out = a_a_ext + a_d_inv;
	wire a_bigger_uneq = unsigned_ == a_a_ext[31];
	wire a_bigger = (a_a_ext[31] == a_d_ext[31] ? ~adder_out[31] : a_bigger_uneq);
	wire pick_a = take_max == a_bigger;
	wire [31:0] _arith_out_T = (pick_a ? cam_a_0_bits_data : cam_d_0_data);
	wire [31:0] arith_out = (adder ? adder_out : _arith_out_T);
	wire [31:0] amo_data = (cam_a_0_bits_opcode[0] ? logic_out : arith_out);
	wire a_allow = ~cam_abusy_0 & (a_isSupported | cam_free_0);
	reg [3:0] beatsLeft;
	wire idle = beatsLeft == 4'h0;
	wire source_i_valid = auto_in_a_valid & a_allow;
	wire [1:0] _readys_T = {source_i_valid, cam_amo_0};
	wire [2:0] _readys_T_1 = {_readys_T, 1'h0};
	wire [1:0] _readys_T_3 = _readys_T | _readys_T_1[1:0];
	wire [2:0] _readys_T_5 = {_readys_T_3, 1'h0};
	wire [1:0] _readys_T_7 = ~_readys_T_5[1:0];
	wire readys_1 = _readys_T_7[1];
	reg state_1;
	wire allowed_1 = (idle ? readys_1 : state_1);
	wire out_1_ready = auto_out_a_ready & allowed_1;
	wire _T = ~a_isSupported;
	wire [2:0] source_i_bits_opcode = (~a_isSupported ? 3'h4 : auto_in_a_bits_opcode);
	wire [2:0] source_i_bits_param = (~a_isSupported ? 3'h0 : auto_in_a_bits_param);
	wire source_c_bits_a_corrupt = cam_a_0_bits_corrupt | cam_d_0_corrupt;
	wire source_c_bits_a_mask_sizeOH_shiftAmount = cam_a_0_bits_size[0];
	wire [1:0] _source_c_bits_a_mask_sizeOH_T_1 = 2'h1 << source_c_bits_a_mask_sizeOH_shiftAmount;
	wire [1:0] source_c_bits_a_mask_sizeOH = _source_c_bits_a_mask_sizeOH_T_1 | 2'h1;
	wire _source_c_bits_a_mask_T = cam_a_0_bits_size >= 3'h2;
	wire source_c_bits_a_mask_size = source_c_bits_a_mask_sizeOH[1];
	wire source_c_bits_a_mask_bit = cam_a_0_bits_address[1];
	wire source_c_bits_a_mask_nbit = ~source_c_bits_a_mask_bit;
	wire source_c_bits_a_mask_acc = _source_c_bits_a_mask_T | (source_c_bits_a_mask_size & source_c_bits_a_mask_nbit);
	wire source_c_bits_a_mask_acc_1 = _source_c_bits_a_mask_T | (source_c_bits_a_mask_size & source_c_bits_a_mask_bit);
	wire source_c_bits_a_mask_size_1 = source_c_bits_a_mask_sizeOH[0];
	wire source_c_bits_a_mask_bit_1 = cam_a_0_bits_address[0];
	wire source_c_bits_a_mask_nbit_1 = ~source_c_bits_a_mask_bit_1;
	wire source_c_bits_a_mask_eq_2 = source_c_bits_a_mask_nbit & source_c_bits_a_mask_nbit_1;
	wire source_c_bits_a_mask_acc_2 = source_c_bits_a_mask_acc | (source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_2);
	wire source_c_bits_a_mask_eq_3 = source_c_bits_a_mask_nbit & source_c_bits_a_mask_bit_1;
	wire source_c_bits_a_mask_acc_3 = source_c_bits_a_mask_acc | (source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_3);
	wire source_c_bits_a_mask_eq_4 = source_c_bits_a_mask_bit & source_c_bits_a_mask_nbit_1;
	wire source_c_bits_a_mask_acc_4 = source_c_bits_a_mask_acc_1 | (source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_4);
	wire source_c_bits_a_mask_eq_5 = source_c_bits_a_mask_bit & source_c_bits_a_mask_bit_1;
	wire source_c_bits_a_mask_acc_5 = source_c_bits_a_mask_acc_1 | (source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_5);
	wire [3:0] source_c_bits_a_mask = {source_c_bits_a_mask_acc_5, source_c_bits_a_mask_acc_4, source_c_bits_a_mask_acc_3, source_c_bits_a_mask_acc_2};
	wire [12:0] _decode_T_1 = 13'h003f << auto_in_a_bits_size;
	wire [5:0] _decode_T_3 = ~_decode_T_1[5:0];
	wire [3:0] decode = _decode_T_3[5:2];
	wire opdata = ~auto_in_a_bits_opcode[2];
	wire latch = idle & auto_out_a_ready;
	wire readys_0 = _readys_T_7[0];
	wire earlyWinner_0 = readys_0 & cam_amo_0;
	wire earlyWinner_1 = readys_1 & source_i_valid;
	wire _prefixOR_T = earlyWinner_0 | earlyWinner_1;
	wire _T_10 = ~reset;
	wire _T_12 = cam_amo_0 | source_i_valid;
	wire _T_13 = ~(cam_amo_0 | source_i_valid);
	reg state_0;
	wire muxStateEarly_0 = (idle ? earlyWinner_0 : state_0);
	wire muxStateEarly_1 = (idle ? earlyWinner_1 : state_1);
	wire _sink_ACancel_earlyValid_T_3 = (state_0 & cam_amo_0) | (state_1 & source_i_valid);
	wire sink_ACancel_earlyValid = (idle ? _T_12 : _sink_ACancel_earlyValid_T_3);
	wire _beatsLeft_T_2 = auto_out_a_ready & sink_ACancel_earlyValid;
	wire [3:0] _GEN_40 = {3'd0, _beatsLeft_T_2};
	wire [3:0] _beatsLeft_T_4 = beatsLeft - _GEN_40;
	wire allowed_0 = (idle ? readys_0 : state_0);
	wire out_ready = auto_out_a_ready & allowed_0;
	wire [31:0] _T_29 = (muxStateEarly_0 ? amo_data : 32'h00000000);
	wire [31:0] _T_30 = (muxStateEarly_1 ? auto_in_a_bits_data : 32'h00000000);
	wire [3:0] _T_32 = (muxStateEarly_0 ? source_c_bits_a_mask : 4'h0);
	wire [3:0] _T_33 = (muxStateEarly_1 ? auto_in_a_bits_mask : 4'h0);
	wire [30:0] _T_35 = (muxStateEarly_0 ? cam_a_0_bits_address : 31'h00000000);
	wire [30:0] _T_36 = (muxStateEarly_1 ? auto_in_a_bits_address : 31'h00000000);
	wire [2:0] _T_38 = (muxStateEarly_0 ? cam_a_0_bits_source : 3'h0);
	wire [2:0] _T_39 = (muxStateEarly_1 ? auto_in_a_bits_source : 3'h0);
	wire [2:0] _T_41 = (muxStateEarly_0 ? cam_a_0_bits_size : 3'h0);
	wire [2:0] _T_42 = (muxStateEarly_1 ? auto_in_a_bits_size : 3'h0);
	wire _T_50 = out_1_ready & source_i_valid;
	wire [2:0] _GEN_41 = {1'd0, auto_in_a_bits_param[1:0]};
	wire [3:0] _cam_a_0_lut_T_2 = (3'h1 == _GEN_41 ? 4'he : 4'h8);
	wire [1:0] _GEN_12 = (cam_free_0 ? 2'h3 : cam_s_0_state);
	wire [1:0] _GEN_23 = (_T_50 & _T ? _GEN_12 : cam_s_0_state);
	wire _T_53 = out_ready & cam_amo_0;
	wire [1:0] _GEN_24 = (cam_amo_0 ? 2'h1 : _GEN_23);
	wire [1:0] _GEN_25 = (_T_53 ? _GEN_24 : _GEN_23);
	reg [3:0] d_first_counter;
	wire d_first = d_first_counter == 4'h0;
	wire d_ackd = auto_out_d_bits_opcode == 3'h1;
	wire d_cam_sel_raw_0 = cam_a_0_bits_source == auto_out_d_bits_source;
	wire d_cam_sel_match_0 = d_cam_sel_raw_0 & cam_dmatch_0;
	wire d_drop = (d_first & d_ackd) & d_cam_sel_match_0;
	wire bundleOut_0_d_ready = auto_in_d_ready | d_drop;
	wire _d_first_T = bundleOut_0_d_ready & auto_out_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << auto_out_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = auto_out_d_bits_opcode[0];
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_ack = auto_out_d_bits_opcode == 3'h0;
	wire d_replace = (d_first & d_ack) & d_cam_sel_match_0;
	TLMonitor_7 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	assign auto_in_a_ready = out_1_ready & a_allow;
	assign auto_in_d_valid = auto_out_d_valid & ~d_drop;
	assign auto_in_d_bits_opcode = (d_replace ? 3'h1 : auto_out_d_bits_opcode);
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = (d_replace ? cam_d_0_denied | auto_out_d_bits_denied : auto_out_d_bits_denied);
	assign auto_in_d_bits_data = (d_replace ? cam_d_0_data : auto_out_d_bits_data);
	assign auto_in_d_bits_corrupt = (d_replace ? cam_d_0_corrupt | auto_out_d_bits_denied : auto_out_d_bits_corrupt);
	assign auto_out_a_valid = (idle ? _T_12 : _sink_ACancel_earlyValid_T_3);
	assign auto_out_a_bits_opcode = (muxStateEarly_1 ? source_i_bits_opcode : 3'h0);
	assign auto_out_a_bits_param = (muxStateEarly_1 ? source_i_bits_param : 3'h0);
	assign auto_out_a_bits_size = _T_41 | _T_42;
	assign auto_out_a_bits_source = _T_38 | _T_39;
	assign auto_out_a_bits_address = _T_35 | _T_36;
	assign auto_out_a_bits_mask = _T_32 | _T_33;
	assign auto_out_a_bits_data = _T_29 | _T_30;
	assign auto_out_a_bits_corrupt = (muxStateEarly_0 & source_c_bits_a_corrupt) | (muxStateEarly_1 & auto_in_a_bits_corrupt);
	assign auto_out_d_ready = auto_in_d_ready | d_drop;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = out_1_ready & a_allow;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid & ~d_drop;
	assign monitor_io_in_d_bits_opcode = (d_replace ? 3'h1 : auto_out_d_bits_opcode);
	assign monitor_io_in_d_bits_param = auto_out_d_bits_param;
	assign monitor_io_in_d_bits_size = auto_out_d_bits_size;
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source;
	assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink;
	assign monitor_io_in_d_bits_denied = (d_replace ? cam_d_0_denied | auto_out_d_bits_denied : auto_out_d_bits_denied);
	assign monitor_io_in_d_bits_corrupt = (d_replace ? cam_d_0_corrupt | auto_out_d_bits_denied : auto_out_d_bits_corrupt);
	always @(posedge clock) begin
		if (reset)
			cam_s_0_state <= 2'h0;
		else if (_d_first_T & d_first) begin
			if (d_cam_sel_match_0) begin
				if (d_ackd)
					cam_s_0_state <= 2'h2;
				else
					cam_s_0_state <= 2'h0;
			end
			else
				cam_s_0_state <= _GEN_25;
		end
		else
			cam_s_0_state <= _GEN_25;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_opcode <= auto_in_a_bits_opcode;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_param <= auto_in_a_bits_param;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_size <= auto_in_a_bits_size;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_source <= auto_in_a_bits_source;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_address <= auto_in_a_bits_address;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_mask <= auto_in_a_bits_mask;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_data <= auto_in_a_bits_data;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_corrupt <= auto_in_a_bits_corrupt;
		if (_T_50 & _T)
			if (cam_free_0)
				if (3'h3 == _GEN_41)
					cam_a_0_lut <= 4'hc;
				else if (3'h0 == _GEN_41)
					cam_a_0_lut <= 4'h6;
				else
					cam_a_0_lut <= _cam_a_0_lut_T_2;
		if (_d_first_T & d_first)
			if (d_cam_sel_match_0 & d_ackd)
				cam_d_0_data <= auto_out_d_bits_data;
		if (_d_first_T & d_first)
			if (d_cam_sel_match_0 & d_ackd)
				cam_d_0_denied <= auto_out_d_bits_denied;
		if (_d_first_T & d_first)
			if (d_cam_sel_match_0 & d_ackd)
				cam_d_0_corrupt <= auto_out_d_bits_corrupt;
		if (reset)
			beatsLeft <= 4'h0;
		else if (latch) begin
			if (earlyWinner_1) begin
				if (opdata)
					beatsLeft <= decode;
				else
					beatsLeft <= 4'h0;
			end
			else
				beatsLeft <= 4'h0;
		end
		else
			beatsLeft <= _beatsLeft_T_4;
		if (reset)
			state_1 <= 1'h0;
		else if (idle)
			state_1 <= earlyWinner_1;
		if (reset)
			state_0 <= 1'h0;
		else if (idle)
			state_0 <= earlyWinner_0;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
	end
endmodule
module TLMonitor_8 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [30:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [30:0] _GEN_71 = {25'd0, is_aligned_mask};
	wire [30:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 31'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [30:0] _T_56 = io_in_a_bits_address ^ 31'h00004000;
	wire [31:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [31:0] _T_59 = $signed(_T_57) & -32'sh00001000;
	wire _T_60 = $signed(_T_59) == 32'sh00000000;
	wire [30:0] _T_61 = io_in_a_bits_address ^ 31'h00020000;
	wire [31:0] _T_62 = {1'b0, $signed(_T_61)};
	wire [31:0] _T_64 = $signed(_T_62) & -32'sh00010000;
	wire _T_65 = $signed(_T_64) == 32'sh00000000;
	wire [30:0] _T_66 = io_in_a_bits_address ^ 31'h10000000;
	wire [31:0] _T_67 = {1'b0, $signed(_T_66)};
	wire [31:0] _T_69 = $signed(_T_67) & -32'sh00001000;
	wire _T_70 = $signed(_T_69) == 32'sh00000000;
	wire [30:0] _T_71 = io_in_a_bits_address ^ 31'h54000000;
	wire [31:0] _T_72 = {1'b0, $signed(_T_71)};
	wire [31:0] _T_74 = $signed(_T_72) & -32'sh00001000;
	wire _T_75 = $signed(_T_74) == 32'sh00000000;
	wire _T_78 = ((_T_60 | _T_65) | _T_70) | _T_75;
	wire _T_128 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_132 = ~io_in_a_bits_mask;
	wire _T_133 = _T_132 == 4'h0;
	wire _T_137 = ~io_in_a_bits_corrupt;
	wire _T_141 = io_in_a_bits_opcode == 3'h7;
	wire _T_231 = io_in_a_bits_param != 3'h0;
	wire _T_244 = io_in_a_bits_opcode == 3'h4;
	wire _T_261 = io_in_a_bits_size <= 3'h6;
	wire _T_287 = _T_261 & _T_78;
	wire _T_298 = io_in_a_bits_param == 3'h0;
	wire _T_302 = io_in_a_bits_mask == mask;
	wire _T_310 = io_in_a_bits_opcode == 3'h0;
	wire _T_343 = (_T_60 | _T_70) | _T_75;
	wire _T_344 = _T_261 & _T_343;
	wire _T_354 = source_ok & _T_344;
	wire _T_372 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_430 = ~mask;
	wire [3:0] _T_431 = io_in_a_bits_mask & _T_430;
	wire _T_432 = _T_431 == 4'h0;
	wire _T_436 = io_in_a_bits_opcode == 3'h2;
	wire _T_450 = io_in_a_bits_size <= 3'h2;
	wire _T_470 = _T_450 & _T_343;
	wire _T_480 = source_ok & _T_470;
	wire _T_490 = io_in_a_bits_param <= 3'h4;
	wire _T_498 = io_in_a_bits_opcode == 3'h3;
	wire _T_552 = io_in_a_bits_param <= 3'h3;
	wire _T_560 = io_in_a_bits_opcode == 3'h5;
	wire _T_609 = io_in_a_bits_param <= 3'h1;
	wire _T_621 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_625 = io_in_d_bits_opcode == 3'h6;
	wire _T_629 = io_in_d_bits_size >= 3'h2;
	wire _T_633 = io_in_d_bits_param == 2'h0;
	wire _T_637 = ~io_in_d_bits_corrupt;
	wire _T_641 = ~io_in_d_bits_denied;
	wire _T_645 = io_in_d_bits_opcode == 3'h4;
	wire _T_656 = io_in_d_bits_param <= 2'h2;
	wire _T_660 = io_in_d_bits_param != 2'h2;
	wire _T_673 = io_in_d_bits_opcode == 3'h5;
	wire _T_693 = _T_641 | io_in_d_bits_corrupt;
	wire _T_702 = io_in_d_bits_opcode == 3'h0;
	wire _T_719 = io_in_d_bits_opcode == 3'h1;
	wire _T_737 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [30:0] address;
	wire _T_767 = io_in_a_valid & ~a_first;
	wire _T_768 = io_in_a_bits_opcode == opcode;
	wire _T_772 = io_in_a_bits_param == param;
	wire _T_776 = io_in_a_bits_size == size;
	wire _T_780 = io_in_a_bits_source == source;
	wire _T_784 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_791 = io_in_d_valid & ~d_first;
	wire _T_792 = io_in_d_bits_opcode == opcode_1;
	wire _T_796 = io_in_d_bits_param == param_1;
	wire _T_800 = io_in_d_bits_size == size_1;
	wire _T_804 = io_in_d_bits_source == source_1;
	wire _T_808 = io_in_d_bits_sink == sink;
	wire _T_812 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_818 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire [7:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire _T_821 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_823 = inflight >> io_in_a_bits_source;
	wire _T_825 = ~_T_823[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_829 = io_in_d_valid & d_first_1;
	wire _T_831 = ~_T_625;
	wire _T_832 = (io_in_d_valid & d_first_1) & ~_T_625;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [7:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_625 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_831 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_831 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_818 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_842 = inflight >> io_in_d_bits_source;
	wire _T_844 = _T_842[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_849 = io_in_d_bits_opcode == _GEN_40;
	wire _T_850 = (io_in_d_bits_opcode == _GEN_32) | _T_849;
	wire _T_854 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_861 = io_in_d_bits_opcode == _GEN_56;
	wire _T_862 = (io_in_d_bits_opcode == _GEN_48) | _T_861;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_866 = _GEN_82 == a_size_lookup;
	wire _T_876 = (((_T_829 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_831;
	wire _T_878 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set_wo_ready = _GEN_15[4:0];
	wire [4:0] d_clr_wo_ready = _GEN_21[4:0];
	wire _T_885 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_894 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_920 = (io_in_d_valid & d_first_2) & _T_625;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_625 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_625 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_928 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_938 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_963 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLBuffer_2 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [30:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [30:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [30:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire bundleOut_0_a_q_clock;
	wire bundleOut_0_a_q_reset;
	wire bundleOut_0_a_q_io_enq_ready;
	wire bundleOut_0_a_q_io_enq_valid;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_param;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_size;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_source;
	wire [30:0] bundleOut_0_a_q_io_enq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_data;
	wire bundleOut_0_a_q_io_enq_bits_corrupt;
	wire bundleOut_0_a_q_io_deq_ready;
	wire bundleOut_0_a_q_io_deq_valid;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_param;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_size;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_source;
	wire [30:0] bundleOut_0_a_q_io_deq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_data;
	wire bundleOut_0_a_q_io_deq_bits_corrupt;
	wire bundleIn_0_d_q_clock;
	wire bundleIn_0_d_q_reset;
	wire bundleIn_0_d_q_io_enq_ready;
	wire bundleIn_0_d_q_io_enq_valid;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_enq_bits_param;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_size;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_source;
	wire bundleIn_0_d_q_io_enq_bits_sink;
	wire bundleIn_0_d_q_io_enq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_enq_bits_data;
	wire bundleIn_0_d_q_io_enq_bits_corrupt;
	wire bundleIn_0_d_q_io_deq_ready;
	wire bundleIn_0_d_q_io_deq_valid;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_param;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_size;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_source;
	wire bundleIn_0_d_q_io_deq_bits_sink;
	wire bundleIn_0_d_q_io_deq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_deq_bits_data;
	wire bundleIn_0_d_q_io_deq_bits_corrupt;
	TLMonitor_8 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Queue bundleOut_0_a_q(
		.clock(bundleOut_0_a_q_clock),
		.reset(bundleOut_0_a_q_reset),
		.io_enq_ready(bundleOut_0_a_q_io_enq_ready),
		.io_enq_valid(bundleOut_0_a_q_io_enq_valid),
		.io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
		.io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
		.io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
		.io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
		.io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
		.io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleOut_0_a_q_io_deq_ready),
		.io_deq_valid(bundleOut_0_a_q_io_deq_valid),
		.io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
		.io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
		.io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
		.io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
		.io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
		.io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
	);
	Queue_1 bundleIn_0_d_q(
		.clock(bundleIn_0_d_q_clock),
		.reset(bundleIn_0_d_q_reset),
		.io_enq_ready(bundleIn_0_d_q_io_enq_ready),
		.io_enq_valid(bundleIn_0_d_q_io_enq_valid),
		.io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
		.io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
		.io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
		.io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
		.io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
		.io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleIn_0_d_q_io_deq_ready),
		.io_deq_valid(bundleIn_0_d_q_io_deq_valid),
		.io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
		.io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
		.io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
		.io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
		.io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
		.io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data;
	assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid;
	assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode;
	assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param;
	assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size;
	assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source;
	assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address;
	assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask;
	assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data;
	assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt;
	assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign bundleOut_0_a_q_clock = clock;
	assign bundleOut_0_a_q_reset = reset;
	assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid;
	assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param;
	assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size;
	assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source;
	assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address;
	assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask;
	assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data;
	assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready;
	assign bundleIn_0_d_q_clock = clock;
	assign bundleIn_0_d_q_reset = reset;
	assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid;
	assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign bundleIn_0_d_q_io_enq_bits_param = auto_out_d_bits_param;
	assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size;
	assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source;
	assign bundleIn_0_d_q_io_enq_bits_sink = auto_out_d_bits_sink;
	assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied;
	assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data;
	assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt;
	assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready;
endmodule
module TLMonitor_9 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [14:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [14:0] _GEN_71 = {9'd0, is_aligned_mask};
	wire [14:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 15'h0000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [14:0] _T_56 = io_in_a_bits_address ^ 15'h4000;
	wire [15:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [15:0] _T_59 = $signed(_T_57) & -16'sh1000;
	wire _T_60 = $signed(_T_59) == 16'sh0000;
	wire _T_92 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_96 = ~io_in_a_bits_mask;
	wire _T_97 = _T_96 == 4'h0;
	wire _T_101 = ~io_in_a_bits_corrupt;
	wire _T_105 = io_in_a_bits_opcode == 3'h7;
	wire _T_159 = io_in_a_bits_param != 3'h0;
	wire _T_172 = io_in_a_bits_opcode == 3'h4;
	wire _T_189 = io_in_a_bits_size <= 3'h6;
	wire _T_197 = _T_189 & _T_60;
	wire _T_208 = io_in_a_bits_param == 3'h0;
	wire _T_212 = io_in_a_bits_mask == mask;
	wire _T_220 = io_in_a_bits_opcode == 3'h0;
	wire _T_244 = source_ok & _T_197;
	wire _T_262 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_300 = ~mask;
	wire [3:0] _T_301 = io_in_a_bits_mask & _T_300;
	wire _T_302 = _T_301 == 4'h0;
	wire _T_306 = io_in_a_bits_opcode == 3'h2;
	wire _T_337 = io_in_a_bits_param <= 3'h4;
	wire _T_345 = io_in_a_bits_opcode == 3'h3;
	wire _T_376 = io_in_a_bits_param <= 3'h3;
	wire _T_384 = io_in_a_bits_opcode == 3'h5;
	wire _T_415 = io_in_a_bits_param <= 3'h1;
	wire _T_427 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_431 = io_in_d_bits_opcode == 3'h6;
	wire _T_435 = io_in_d_bits_size >= 3'h2;
	wire _T_451 = io_in_d_bits_opcode == 3'h4;
	wire _T_479 = io_in_d_bits_opcode == 3'h5;
	wire _T_508 = io_in_d_bits_opcode == 3'h0;
	wire _T_525 = io_in_d_bits_opcode == 3'h1;
	wire _T_543 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [14:0] address;
	wire _T_573 = io_in_a_valid & ~a_first;
	wire _T_574 = io_in_a_bits_opcode == opcode;
	wire _T_578 = io_in_a_bits_param == param;
	wire _T_582 = io_in_a_bits_size == size;
	wire _T_586 = io_in_a_bits_source == source;
	wire _T_590 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	wire _T_597 = io_in_d_valid & ~d_first;
	wire _T_598 = io_in_d_bits_opcode == opcode_1;
	wire _T_606 = io_in_d_bits_size == size_1;
	wire _T_610 = io_in_d_bits_source == source_1;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_624 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire _T_627 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_629 = inflight >> io_in_a_bits_source;
	wire _T_631 = ~_T_629[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_635 = io_in_d_valid & d_first_1;
	wire _T_637 = ~_T_431;
	wire _T_638 = (io_in_d_valid & d_first_1) & ~_T_431;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_637 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_637 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_624 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_648 = inflight >> io_in_d_bits_source;
	wire _T_650 = _T_648[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_655 = io_in_d_bits_opcode == _GEN_40;
	wire _T_656 = (io_in_d_bits_opcode == _GEN_32) | _T_655;
	wire _T_660 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_667 = io_in_d_bits_opcode == _GEN_56;
	wire _T_668 = (io_in_d_bits_opcode == _GEN_48) | _T_667;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_672 = _GEN_82 == a_size_lookup;
	wire _T_682 = (((_T_635 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_637;
	wire _T_684 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_693 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_719 = (io_in_d_valid & d_first_2) & _T_431;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_431 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_431 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_727 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_737 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_757 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Repeater (
	clock,
	reset,
	io_repeat,
	io_full,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	input io_repeat;
	output wire io_full;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [14:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [14:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire io_deq_bits_corrupt;
	reg full;
	reg [2:0] saved_opcode;
	reg [2:0] saved_param;
	reg [2:0] saved_size;
	reg [2:0] saved_source;
	reg [14:0] saved_address;
	reg [3:0] saved_mask;
	reg saved_corrupt;
	wire _T = io_enq_ready & io_enq_valid;
	wire _GEN_0 = (_T & io_repeat) | full;
	wire _T_2 = io_deq_ready & io_deq_valid;
	assign io_full = full;
	assign io_enq_ready = io_deq_ready & ~full;
	assign io_deq_valid = io_enq_valid | full;
	assign io_deq_bits_opcode = (full ? saved_opcode : io_enq_bits_opcode);
	assign io_deq_bits_param = (full ? saved_param : io_enq_bits_param);
	assign io_deq_bits_size = (full ? saved_size : io_enq_bits_size);
	assign io_deq_bits_source = (full ? saved_source : io_enq_bits_source);
	assign io_deq_bits_address = (full ? saved_address : io_enq_bits_address);
	assign io_deq_bits_mask = (full ? saved_mask : io_enq_bits_mask);
	assign io_deq_bits_corrupt = (full ? saved_corrupt : io_enq_bits_corrupt);
	always @(posedge clock) begin
		if (reset)
			full <= 1'h0;
		else if (_T_2 & ~io_repeat)
			full <= 1'h0;
		else
			full <= _GEN_0;
		if (_T & io_repeat)
			saved_opcode <= io_enq_bits_opcode;
		if (_T & io_repeat)
			saved_param <= io_enq_bits_param;
		if (_T & io_repeat)
			saved_size <= io_enq_bits_size;
		if (_T & io_repeat)
			saved_source <= io_enq_bits_source;
		if (_T & io_repeat)
			saved_address <= io_enq_bits_address;
		if (_T & io_repeat)
			saved_mask <= io_enq_bits_mask;
		if (_T & io_repeat)
			saved_corrupt <= io_enq_bits_corrupt;
	end
endmodule
module TLFragmenter (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [14:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire [7:0] auto_out_a_bits_source;
	output wire [14:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_size;
	input [7:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [14:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire repeater_clock;
	wire repeater_reset;
	wire repeater_io_repeat;
	wire repeater_io_full;
	wire repeater_io_enq_ready;
	wire repeater_io_enq_valid;
	wire [2:0] repeater_io_enq_bits_opcode;
	wire [2:0] repeater_io_enq_bits_param;
	wire [2:0] repeater_io_enq_bits_size;
	wire [2:0] repeater_io_enq_bits_source;
	wire [14:0] repeater_io_enq_bits_address;
	wire [3:0] repeater_io_enq_bits_mask;
	wire repeater_io_enq_bits_corrupt;
	wire repeater_io_deq_ready;
	wire repeater_io_deq_valid;
	wire [2:0] repeater_io_deq_bits_opcode;
	wire [2:0] repeater_io_deq_bits_param;
	wire [2:0] repeater_io_deq_bits_size;
	wire [2:0] repeater_io_deq_bits_source;
	wire [14:0] repeater_io_deq_bits_address;
	wire [3:0] repeater_io_deq_bits_mask;
	wire repeater_io_deq_bits_corrupt;
	reg [3:0] acknum;
	reg [2:0] dOrig;
	reg dToggle;
	wire [3:0] dFragnum = auto_out_d_bits_source[3:0];
	wire dFirst = acknum == 4'h0;
	wire dLast = dFragnum == 4'h0;
	wire [3:0] _dsizeOH_T = 4'h1 << auto_out_d_bits_size;
	wire [2:0] dsizeOH = _dsizeOH_T[2:0];
	wire [4:0] _dsizeOH1_T_1 = 5'h03 << auto_out_d_bits_size;
	wire [1:0] dsizeOH1 = ~_dsizeOH1_T_1[1:0];
	wire dHasData = auto_out_d_bits_opcode[0];
	wire _T_5 = ~reset;
	wire ack_decrement = dHasData | dsizeOH[2];
	wire [5:0] _dFirst_size_T = {dFragnum, 2'h0};
	wire [5:0] _GEN_7 = {4'd0, dsizeOH1};
	wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7;
	wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0};
	wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h01;
	wire [6:0] _dFirst_size_T_4 = {1'h0, _dFirst_size_T_1};
	wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4;
	wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5;
	wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4];
	wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0];
	wire _dFirst_size_T_7 = |dFirst_size_hi;
	wire [3:0] _GEN_8 = {1'd0, dFirst_size_hi};
	wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo;
	wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2];
	wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0];
	wire _dFirst_size_T_9 = |dFirst_size_hi_1;
	wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1;
	wire [2:0] dFirst_size = {_dFirst_size_T_7, _dFirst_size_T_9, _dFirst_size_T_10[1]};
	wire drop = ~dHasData & ~dLast;
	wire bundleOut_0_d_ready = auto_in_d_ready | drop;
	wire _T_7 = bundleOut_0_d_ready & auto_out_d_valid;
	wire [3:0] _GEN_9 = {3'd0, ack_decrement};
	wire [3:0] _acknum_T_1 = acknum - _GEN_9;
	wire [2:0] aFrag = (repeater_io_deq_bits_size > 3'h2 ? 3'h2 : repeater_io_deq_bits_size);
	wire [12:0] _aOrigOH1_T_1 = 13'h003f << repeater_io_deq_bits_size;
	wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0];
	wire [8:0] _aFragOH1_T_1 = 9'h003 << aFrag;
	wire [1:0] aFragOH1 = ~_aFragOH1_T_1[1:0];
	wire aHasData = ~repeater_io_deq_bits_opcode[2];
	reg [3:0] gennum;
	wire aFirst = gennum == 4'h0;
	wire [3:0] _old_gennum1_T_2 = gennum - 4'h1;
	wire [3:0] old_gennum1 = (aFirst ? aOrigOH1[5:2] : _old_gennum1_T_2);
	wire [3:0] _new_gennum_T = ~old_gennum1;
	wire [3:0] new_gennum = ~_new_gennum_T;
	reg aToggle_r;
	wire _GEN_5 = (aFirst ? dToggle : aToggle_r);
	wire aToggle = ~_GEN_5;
	wire bundleOut_0_a_valid = repeater_io_deq_valid;
	wire _T_8 = auto_out_a_ready & bundleOut_0_a_valid;
	wire _repeater_io_repeat_T = ~aHasData;
	wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 2'h0};
	wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1;
	wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1;
	wire [5:0] _GEN_10 = {4'd0, aFragOH1};
	wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10;
	wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h03;
	wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4;
	wire [14:0] _GEN_11 = {9'd0, _bundleOut_0_a_bits_address_T_5};
	wire [3:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source, aToggle};
	wire _T_9 = ~repeater_io_full;
	TLMonitor_9 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	Repeater repeater(
		.clock(repeater_clock),
		.reset(repeater_reset),
		.io_repeat(repeater_io_repeat),
		.io_full(repeater_io_full),
		.io_enq_ready(repeater_io_enq_ready),
		.io_enq_valid(repeater_io_enq_valid),
		.io_enq_bits_opcode(repeater_io_enq_bits_opcode),
		.io_enq_bits_param(repeater_io_enq_bits_param),
		.io_enq_bits_size(repeater_io_enq_bits_size),
		.io_enq_bits_source(repeater_io_enq_bits_source),
		.io_enq_bits_address(repeater_io_enq_bits_address),
		.io_enq_bits_mask(repeater_io_enq_bits_mask),
		.io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
		.io_deq_ready(repeater_io_deq_ready),
		.io_deq_valid(repeater_io_deq_valid),
		.io_deq_bits_opcode(repeater_io_deq_bits_opcode),
		.io_deq_bits_param(repeater_io_deq_bits_param),
		.io_deq_bits_size(repeater_io_deq_bits_size),
		.io_deq_bits_source(repeater_io_deq_bits_source),
		.io_deq_bits_address(repeater_io_deq_bits_address),
		.io_deq_bits_mask(repeater_io_deq_bits_mask),
		.io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = repeater_io_enq_ready;
	assign auto_in_d_valid = auto_out_d_valid & ~drop;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign auto_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_out_a_valid = repeater_io_deq_valid;
	assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode;
	assign auto_out_a_bits_param = repeater_io_deq_bits_param;
	assign auto_out_a_bits_size = aFrag[1:0];
	assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi, new_gennum};
	assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11;
	assign auto_out_a_bits_mask = (repeater_io_full ? 4'hf : auto_in_a_bits_mask);
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready | drop;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = repeater_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid & ~drop;
	assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_io_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign repeater_clock = clock;
	assign repeater_reset = reset;
	assign repeater_io_repeat = ~aHasData & (new_gennum != 4'h0);
	assign repeater_io_enq_valid = auto_in_a_valid;
	assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign repeater_io_enq_bits_param = auto_in_a_bits_param;
	assign repeater_io_enq_bits_size = auto_in_a_bits_size;
	assign repeater_io_enq_bits_source = auto_in_a_bits_source;
	assign repeater_io_enq_bits_address = auto_in_a_bits_address;
	assign repeater_io_enq_bits_mask = auto_in_a_bits_mask;
	assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign repeater_io_deq_ready = auto_out_a_ready;
	always @(posedge clock) begin
		if (reset)
			acknum <= 4'h0;
		else if (_T_7)
			if (dFirst)
				acknum <= dFragnum;
			else
				acknum <= _acknum_T_1;
		if (_T_7)
			if (dFirst)
				dOrig <= dFirst_size;
		if (reset)
			dToggle <= 1'h0;
		else if (_T_7)
			if (dFirst)
				dToggle <= auto_out_d_bits_source[4];
		if (reset)
			gennum <= 4'h0;
		else if (_T_8)
			gennum <= new_gennum;
		if (aFirst)
			aToggle_r <= dToggle;
	end
endmodule
module TLBuffer_3 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [14:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [14:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module TLInterconnectCoupler_5 (
	clock,
	reset,
	auto_buffer_in_a_ready,
	auto_buffer_in_a_valid,
	auto_buffer_in_a_bits_opcode,
	auto_buffer_in_a_bits_param,
	auto_buffer_in_a_bits_size,
	auto_buffer_in_a_bits_source,
	auto_buffer_in_a_bits_address,
	auto_buffer_in_a_bits_mask,
	auto_buffer_in_a_bits_data,
	auto_buffer_in_a_bits_corrupt,
	auto_buffer_in_d_ready,
	auto_buffer_in_d_valid,
	auto_buffer_in_d_bits_opcode,
	auto_buffer_in_d_bits_size,
	auto_buffer_in_d_bits_source,
	auto_buffer_in_d_bits_data,
	auto_fragmenter_out_a_ready,
	auto_fragmenter_out_a_valid,
	auto_fragmenter_out_a_bits_opcode,
	auto_fragmenter_out_a_bits_param,
	auto_fragmenter_out_a_bits_size,
	auto_fragmenter_out_a_bits_source,
	auto_fragmenter_out_a_bits_address,
	auto_fragmenter_out_a_bits_mask,
	auto_fragmenter_out_a_bits_data,
	auto_fragmenter_out_a_bits_corrupt,
	auto_fragmenter_out_d_ready,
	auto_fragmenter_out_d_valid,
	auto_fragmenter_out_d_bits_opcode,
	auto_fragmenter_out_d_bits_size,
	auto_fragmenter_out_d_bits_source,
	auto_fragmenter_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_buffer_in_a_ready;
	input auto_buffer_in_a_valid;
	input [2:0] auto_buffer_in_a_bits_opcode;
	input [2:0] auto_buffer_in_a_bits_param;
	input [2:0] auto_buffer_in_a_bits_size;
	input [2:0] auto_buffer_in_a_bits_source;
	input [14:0] auto_buffer_in_a_bits_address;
	input [3:0] auto_buffer_in_a_bits_mask;
	input [31:0] auto_buffer_in_a_bits_data;
	input auto_buffer_in_a_bits_corrupt;
	input auto_buffer_in_d_ready;
	output wire auto_buffer_in_d_valid;
	output wire [2:0] auto_buffer_in_d_bits_opcode;
	output wire [2:0] auto_buffer_in_d_bits_size;
	output wire [2:0] auto_buffer_in_d_bits_source;
	output wire [31:0] auto_buffer_in_d_bits_data;
	input auto_fragmenter_out_a_ready;
	output wire auto_fragmenter_out_a_valid;
	output wire [2:0] auto_fragmenter_out_a_bits_opcode;
	output wire [2:0] auto_fragmenter_out_a_bits_param;
	output wire [1:0] auto_fragmenter_out_a_bits_size;
	output wire [7:0] auto_fragmenter_out_a_bits_source;
	output wire [14:0] auto_fragmenter_out_a_bits_address;
	output wire [3:0] auto_fragmenter_out_a_bits_mask;
	output wire [31:0] auto_fragmenter_out_a_bits_data;
	output wire auto_fragmenter_out_a_bits_corrupt;
	output wire auto_fragmenter_out_d_ready;
	input auto_fragmenter_out_d_valid;
	input [2:0] auto_fragmenter_out_d_bits_opcode;
	input [1:0] auto_fragmenter_out_d_bits_size;
	input [7:0] auto_fragmenter_out_d_bits_source;
	input [31:0] auto_fragmenter_out_d_bits_data;
	wire fragmenter_clock;
	wire fragmenter_reset;
	wire fragmenter_auto_in_a_ready;
	wire fragmenter_auto_in_a_valid;
	wire [2:0] fragmenter_auto_in_a_bits_opcode;
	wire [2:0] fragmenter_auto_in_a_bits_param;
	wire [2:0] fragmenter_auto_in_a_bits_size;
	wire [2:0] fragmenter_auto_in_a_bits_source;
	wire [14:0] fragmenter_auto_in_a_bits_address;
	wire [3:0] fragmenter_auto_in_a_bits_mask;
	wire [31:0] fragmenter_auto_in_a_bits_data;
	wire fragmenter_auto_in_a_bits_corrupt;
	wire fragmenter_auto_in_d_ready;
	wire fragmenter_auto_in_d_valid;
	wire [2:0] fragmenter_auto_in_d_bits_opcode;
	wire [2:0] fragmenter_auto_in_d_bits_size;
	wire [2:0] fragmenter_auto_in_d_bits_source;
	wire [31:0] fragmenter_auto_in_d_bits_data;
	wire fragmenter_auto_out_a_ready;
	wire fragmenter_auto_out_a_valid;
	wire [2:0] fragmenter_auto_out_a_bits_opcode;
	wire [2:0] fragmenter_auto_out_a_bits_param;
	wire [1:0] fragmenter_auto_out_a_bits_size;
	wire [7:0] fragmenter_auto_out_a_bits_source;
	wire [14:0] fragmenter_auto_out_a_bits_address;
	wire [3:0] fragmenter_auto_out_a_bits_mask;
	wire [31:0] fragmenter_auto_out_a_bits_data;
	wire fragmenter_auto_out_a_bits_corrupt;
	wire fragmenter_auto_out_d_ready;
	wire fragmenter_auto_out_d_valid;
	wire [2:0] fragmenter_auto_out_d_bits_opcode;
	wire [1:0] fragmenter_auto_out_d_bits_size;
	wire [7:0] fragmenter_auto_out_d_bits_source;
	wire [31:0] fragmenter_auto_out_d_bits_data;
	wire buffer_auto_in_a_ready;
	wire buffer_auto_in_a_valid;
	wire [2:0] buffer_auto_in_a_bits_opcode;
	wire [2:0] buffer_auto_in_a_bits_param;
	wire [2:0] buffer_auto_in_a_bits_size;
	wire [2:0] buffer_auto_in_a_bits_source;
	wire [14:0] buffer_auto_in_a_bits_address;
	wire [3:0] buffer_auto_in_a_bits_mask;
	wire [31:0] buffer_auto_in_a_bits_data;
	wire buffer_auto_in_a_bits_corrupt;
	wire buffer_auto_in_d_ready;
	wire buffer_auto_in_d_valid;
	wire [2:0] buffer_auto_in_d_bits_opcode;
	wire [2:0] buffer_auto_in_d_bits_size;
	wire [2:0] buffer_auto_in_d_bits_source;
	wire [31:0] buffer_auto_in_d_bits_data;
	wire buffer_auto_out_a_ready;
	wire buffer_auto_out_a_valid;
	wire [2:0] buffer_auto_out_a_bits_opcode;
	wire [2:0] buffer_auto_out_a_bits_param;
	wire [2:0] buffer_auto_out_a_bits_size;
	wire [2:0] buffer_auto_out_a_bits_source;
	wire [14:0] buffer_auto_out_a_bits_address;
	wire [3:0] buffer_auto_out_a_bits_mask;
	wire [31:0] buffer_auto_out_a_bits_data;
	wire buffer_auto_out_a_bits_corrupt;
	wire buffer_auto_out_d_ready;
	wire buffer_auto_out_d_valid;
	wire [2:0] buffer_auto_out_d_bits_opcode;
	wire [2:0] buffer_auto_out_d_bits_size;
	wire [2:0] buffer_auto_out_d_bits_source;
	wire [31:0] buffer_auto_out_d_bits_data;
	TLFragmenter fragmenter(
		.clock(fragmenter_clock),
		.reset(fragmenter_reset),
		.auto_in_a_ready(fragmenter_auto_in_a_ready),
		.auto_in_a_valid(fragmenter_auto_in_a_valid),
		.auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
		.auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
		.auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
		.auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
		.auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
		.auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
		.auto_in_d_ready(fragmenter_auto_in_d_ready),
		.auto_in_d_valid(fragmenter_auto_in_d_valid),
		.auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
		.auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
		.auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
		.auto_out_a_ready(fragmenter_auto_out_a_ready),
		.auto_out_a_valid(fragmenter_auto_out_a_valid),
		.auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
		.auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
		.auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
		.auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
		.auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
		.auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
		.auto_out_d_ready(fragmenter_auto_out_d_ready),
		.auto_out_d_valid(fragmenter_auto_out_d_valid),
		.auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
		.auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
		.auto_out_d_bits_data(fragmenter_auto_out_d_bits_data)
	);
	TLBuffer_3 buffer(
		.auto_in_a_ready(buffer_auto_in_a_ready),
		.auto_in_a_valid(buffer_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_auto_in_d_ready),
		.auto_in_d_valid(buffer_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(buffer_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_auto_in_d_bits_source),
		.auto_in_d_bits_data(buffer_auto_in_d_bits_data),
		.auto_out_a_ready(buffer_auto_out_a_ready),
		.auto_out_a_valid(buffer_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_auto_out_d_ready),
		.auto_out_d_valid(buffer_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(buffer_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_auto_out_d_bits_source),
		.auto_out_d_bits_data(buffer_auto_out_d_bits_data)
	);
	assign auto_buffer_in_a_ready = buffer_auto_in_a_ready;
	assign auto_buffer_in_d_valid = buffer_auto_in_d_valid;
	assign auto_buffer_in_d_bits_opcode = buffer_auto_in_d_bits_opcode;
	assign auto_buffer_in_d_bits_size = buffer_auto_in_d_bits_size;
	assign auto_buffer_in_d_bits_source = buffer_auto_in_d_bits_source;
	assign auto_buffer_in_d_bits_data = buffer_auto_in_d_bits_data;
	assign auto_fragmenter_out_a_valid = fragmenter_auto_out_a_valid;
	assign auto_fragmenter_out_a_bits_opcode = fragmenter_auto_out_a_bits_opcode;
	assign auto_fragmenter_out_a_bits_param = fragmenter_auto_out_a_bits_param;
	assign auto_fragmenter_out_a_bits_size = fragmenter_auto_out_a_bits_size;
	assign auto_fragmenter_out_a_bits_source = fragmenter_auto_out_a_bits_source;
	assign auto_fragmenter_out_a_bits_address = fragmenter_auto_out_a_bits_address;
	assign auto_fragmenter_out_a_bits_mask = fragmenter_auto_out_a_bits_mask;
	assign auto_fragmenter_out_a_bits_data = fragmenter_auto_out_a_bits_data;
	assign auto_fragmenter_out_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt;
	assign auto_fragmenter_out_d_ready = fragmenter_auto_out_d_ready;
	assign fragmenter_clock = clock;
	assign fragmenter_reset = reset;
	assign fragmenter_auto_in_a_valid = buffer_auto_out_a_valid;
	assign fragmenter_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode;
	assign fragmenter_auto_in_a_bits_param = buffer_auto_out_a_bits_param;
	assign fragmenter_auto_in_a_bits_size = buffer_auto_out_a_bits_size;
	assign fragmenter_auto_in_a_bits_source = buffer_auto_out_a_bits_source;
	assign fragmenter_auto_in_a_bits_address = buffer_auto_out_a_bits_address;
	assign fragmenter_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask;
	assign fragmenter_auto_in_a_bits_data = buffer_auto_out_a_bits_data;
	assign fragmenter_auto_in_a_bits_corrupt = buffer_auto_out_a_bits_corrupt;
	assign fragmenter_auto_in_d_ready = buffer_auto_out_d_ready;
	assign fragmenter_auto_out_a_ready = auto_fragmenter_out_a_ready;
	assign fragmenter_auto_out_d_valid = auto_fragmenter_out_d_valid;
	assign fragmenter_auto_out_d_bits_opcode = auto_fragmenter_out_d_bits_opcode;
	assign fragmenter_auto_out_d_bits_size = auto_fragmenter_out_d_bits_size;
	assign fragmenter_auto_out_d_bits_source = auto_fragmenter_out_d_bits_source;
	assign fragmenter_auto_out_d_bits_data = auto_fragmenter_out_d_bits_data;
	assign buffer_auto_in_a_valid = auto_buffer_in_a_valid;
	assign buffer_auto_in_a_bits_opcode = auto_buffer_in_a_bits_opcode;
	assign buffer_auto_in_a_bits_param = auto_buffer_in_a_bits_param;
	assign buffer_auto_in_a_bits_size = auto_buffer_in_a_bits_size;
	assign buffer_auto_in_a_bits_source = auto_buffer_in_a_bits_source;
	assign buffer_auto_in_a_bits_address = auto_buffer_in_a_bits_address;
	assign buffer_auto_in_a_bits_mask = auto_buffer_in_a_bits_mask;
	assign buffer_auto_in_a_bits_data = auto_buffer_in_a_bits_data;
	assign buffer_auto_in_a_bits_corrupt = auto_buffer_in_a_bits_corrupt;
	assign buffer_auto_in_d_ready = auto_buffer_in_d_ready;
	assign buffer_auto_out_a_ready = fragmenter_auto_in_a_ready;
	assign buffer_auto_out_d_valid = fragmenter_auto_in_d_valid;
	assign buffer_auto_out_d_bits_opcode = fragmenter_auto_in_d_bits_opcode;
	assign buffer_auto_out_d_bits_size = fragmenter_auto_in_d_bits_size;
	assign buffer_auto_out_d_bits_source = fragmenter_auto_in_d_bits_source;
	assign buffer_auto_out_d_bits_data = fragmenter_auto_in_d_bits_data;
endmodule
module TLSourceShrinker_1 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [28:0] auto_in_a_bits_address;
	input [7:0] auto_in_a_bits_mask;
	input [63:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [63:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [28:0] auto_out_a_bits_address;
	output wire [7:0] auto_out_a_bits_mask;
	output wire [63:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [63:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module TLMonitor_10 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [28:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [28:0] _GEN_71 = {23'd0, is_aligned_mask};
	wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 29'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [28:0] _T_56 = io_in_a_bits_address ^ 29'h00020000;
	wire [29:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [29:0] _T_59 = $signed(_T_57) & -30'sh00010000;
	wire _T_60 = $signed(_T_59) == 30'sh00000000;
	wire [28:0] _T_61 = io_in_a_bits_address ^ 29'h10000000;
	wire [29:0] _T_62 = {1'b0, $signed(_T_61)};
	wire [29:0] _T_64 = $signed(_T_62) & -30'sh00001000;
	wire _T_65 = $signed(_T_64) == 30'sh00000000;
	wire _T_66 = _T_60 | _T_65;
	wire _T_104 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_108 = ~io_in_a_bits_mask;
	wire _T_109 = _T_108 == 4'h0;
	wire _T_113 = ~io_in_a_bits_corrupt;
	wire _T_117 = io_in_a_bits_opcode == 3'h7;
	wire _T_183 = io_in_a_bits_param != 3'h0;
	wire _T_196 = io_in_a_bits_opcode == 3'h4;
	wire _T_213 = io_in_a_bits_size <= 3'h6;
	wire _T_227 = _T_213 & _T_66;
	wire _T_238 = io_in_a_bits_param == 3'h0;
	wire _T_242 = io_in_a_bits_mask == mask;
	wire _T_250 = io_in_a_bits_opcode == 3'h0;
	wire _T_272 = _T_213 & _T_65;
	wire _T_282 = source_ok & _T_272;
	wire _T_300 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_346 = ~mask;
	wire [3:0] _T_347 = io_in_a_bits_mask & _T_346;
	wire _T_348 = _T_347 == 4'h0;
	wire _T_352 = io_in_a_bits_opcode == 3'h2;
	wire _T_389 = io_in_a_bits_param <= 3'h4;
	wire _T_397 = io_in_a_bits_opcode == 3'h3;
	wire _T_434 = io_in_a_bits_param <= 3'h3;
	wire _T_442 = io_in_a_bits_opcode == 3'h5;
	wire _T_479 = io_in_a_bits_param <= 3'h1;
	wire _T_491 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_495 = io_in_d_bits_opcode == 3'h6;
	wire _T_499 = io_in_d_bits_size >= 3'h2;
	wire _T_503 = io_in_d_bits_param == 2'h0;
	wire _T_507 = ~io_in_d_bits_corrupt;
	wire _T_511 = ~io_in_d_bits_denied;
	wire _T_515 = io_in_d_bits_opcode == 3'h4;
	wire _T_526 = io_in_d_bits_param <= 2'h2;
	wire _T_530 = io_in_d_bits_param != 2'h2;
	wire _T_543 = io_in_d_bits_opcode == 3'h5;
	wire _T_563 = _T_511 | io_in_d_bits_corrupt;
	wire _T_572 = io_in_d_bits_opcode == 3'h0;
	wire _T_589 = io_in_d_bits_opcode == 3'h1;
	wire _T_607 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [28:0] address;
	wire _T_637 = io_in_a_valid & ~a_first;
	wire _T_638 = io_in_a_bits_opcode == opcode;
	wire _T_642 = io_in_a_bits_param == param;
	wire _T_646 = io_in_a_bits_size == size;
	wire _T_650 = io_in_a_bits_source == source;
	wire _T_654 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_661 = io_in_d_valid & ~d_first;
	wire _T_662 = io_in_d_bits_opcode == opcode_1;
	wire _T_666 = io_in_d_bits_param == param_1;
	wire _T_670 = io_in_d_bits_size == size_1;
	wire _T_674 = io_in_d_bits_source == source_1;
	wire _T_678 = io_in_d_bits_sink == sink;
	wire _T_682 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_688 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire [7:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire _T_691 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_693 = inflight >> io_in_a_bits_source;
	wire _T_695 = ~_T_693[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_699 = io_in_d_valid & d_first_1;
	wire _T_701 = ~_T_495;
	wire _T_702 = (io_in_d_valid & d_first_1) & ~_T_495;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [7:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_495 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_701 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_701 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_688 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_712 = inflight >> io_in_d_bits_source;
	wire _T_714 = _T_712[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_719 = io_in_d_bits_opcode == _GEN_40;
	wire _T_720 = (io_in_d_bits_opcode == _GEN_32) | _T_719;
	wire _T_724 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_731 = io_in_d_bits_opcode == _GEN_56;
	wire _T_732 = (io_in_d_bits_opcode == _GEN_48) | _T_731;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_736 = _GEN_82 == a_size_lookup;
	wire _T_746 = (((_T_699 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_701;
	wire _T_748 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set_wo_ready = _GEN_15[4:0];
	wire [4:0] d_clr_wo_ready = _GEN_21[4:0];
	wire _T_755 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_764 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_790 = (io_in_d_valid & d_first_2) & _T_495;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_495 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_495 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_798 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_808 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_833 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Repeater_1 (
	clock,
	reset,
	io_repeat,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_sink,
	io_enq_bits_denied,
	io_enq_bits_data,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_sink,
	io_deq_bits_denied,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	input io_repeat;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [1:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input io_enq_bits_sink;
	input io_enq_bits_denied;
	input [63:0] io_enq_bits_data;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [1:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire io_deq_bits_sink;
	output wire io_deq_bits_denied;
	output wire [63:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg full;
	reg [2:0] saved_opcode;
	reg [1:0] saved_param;
	reg [2:0] saved_size;
	reg [2:0] saved_source;
	reg saved_sink;
	reg saved_denied;
	reg [63:0] saved_data;
	reg saved_corrupt;
	wire _T = io_enq_ready & io_enq_valid;
	wire _GEN_0 = (_T & io_repeat) | full;
	wire _T_2 = io_deq_ready & io_deq_valid;
	assign io_enq_ready = io_deq_ready & ~full;
	assign io_deq_valid = io_enq_valid | full;
	assign io_deq_bits_opcode = (full ? saved_opcode : io_enq_bits_opcode);
	assign io_deq_bits_param = (full ? saved_param : io_enq_bits_param);
	assign io_deq_bits_size = (full ? saved_size : io_enq_bits_size);
	assign io_deq_bits_source = (full ? saved_source : io_enq_bits_source);
	assign io_deq_bits_sink = (full ? saved_sink : io_enq_bits_sink);
	assign io_deq_bits_denied = (full ? saved_denied : io_enq_bits_denied);
	assign io_deq_bits_data = (full ? saved_data : io_enq_bits_data);
	assign io_deq_bits_corrupt = (full ? saved_corrupt : io_enq_bits_corrupt);
	always @(posedge clock) begin
		if (reset)
			full <= 1'h0;
		else if (_T_2 & ~io_repeat)
			full <= 1'h0;
		else
			full <= _GEN_0;
		if (_T & io_repeat)
			saved_opcode <= io_enq_bits_opcode;
		if (_T & io_repeat)
			saved_param <= io_enq_bits_param;
		if (_T & io_repeat)
			saved_size <= io_enq_bits_size;
		if (_T & io_repeat)
			saved_source <= io_enq_bits_source;
		if (_T & io_repeat)
			saved_sink <= io_enq_bits_sink;
		if (_T & io_repeat)
			saved_denied <= io_enq_bits_denied;
		if (_T & io_repeat)
			saved_data <= io_enq_bits_data;
		if (_T & io_repeat)
			saved_corrupt <= io_enq_bits_corrupt;
	end
endmodule
module TLWidthWidget_4 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [28:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [28:0] auto_out_a_bits_address;
	output wire [7:0] auto_out_a_bits_mask;
	output wire [63:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [63:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [28:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire repeated_repeater_clock;
	wire repeated_repeater_reset;
	wire repeated_repeater_io_repeat;
	wire repeated_repeater_io_enq_ready;
	wire repeated_repeater_io_enq_valid;
	wire [2:0] repeated_repeater_io_enq_bits_opcode;
	wire [1:0] repeated_repeater_io_enq_bits_param;
	wire [2:0] repeated_repeater_io_enq_bits_size;
	wire [2:0] repeated_repeater_io_enq_bits_source;
	wire repeated_repeater_io_enq_bits_sink;
	wire repeated_repeater_io_enq_bits_denied;
	wire [63:0] repeated_repeater_io_enq_bits_data;
	wire repeated_repeater_io_enq_bits_corrupt;
	wire repeated_repeater_io_deq_ready;
	wire repeated_repeater_io_deq_valid;
	wire [2:0] repeated_repeater_io_deq_bits_opcode;
	wire [1:0] repeated_repeater_io_deq_bits_param;
	wire [2:0] repeated_repeater_io_deq_bits_size;
	wire [2:0] repeated_repeater_io_deq_bits_source;
	wire repeated_repeater_io_deq_bits_sink;
	wire repeated_repeater_io_deq_bits_denied;
	wire [63:0] repeated_repeater_io_deq_bits_data;
	wire repeated_repeater_io_deq_bits_corrupt;
	wire hasData = ~auto_in_a_bits_opcode[2];
	wire [9:0] _limit_T_1 = 10'h007 << auto_in_a_bits_size;
	wire [2:0] _limit_T_3 = ~_limit_T_1[2:0];
	wire limit = _limit_T_3[2];
	reg count;
	wire last = (count == limit) | ~hasData;
	wire enable_0 = ~(|(count & limit));
	reg corrupt_reg;
	wire corrupt_out = auto_in_a_bits_corrupt | corrupt_reg;
	wire _bundleIn_0_a_ready_T = ~last;
	wire bundleIn_0_a_ready = auto_out_a_ready | ~last;
	wire _T = bundleIn_0_a_ready & auto_in_a_valid;
	reg bundleOut_0_a_bits_data_rdata_written_once;
	wire bundleOut_0_a_bits_data_masked_enable_0 = enable_0 | ~bundleOut_0_a_bits_data_rdata_written_once;
	reg [31:0] bundleOut_0_a_bits_data_rdata_0;
	wire [31:0] bundleOut_0_a_bits_data_mdata_0 = (bundleOut_0_a_bits_data_masked_enable_0 ? auto_in_a_bits_data : bundleOut_0_a_bits_data_rdata_0);
	wire _GEN_4 = (_T & _bundleIn_0_a_ready_T) | bundleOut_0_a_bits_data_rdata_written_once;
	wire [1:0] bundleOut_0_a_bits_mask_sizeOH_shiftAmount = auto_in_a_bits_size[1:0];
	wire [3:0] _bundleOut_0_a_bits_mask_sizeOH_T_1 = 4'h1 << bundleOut_0_a_bits_mask_sizeOH_shiftAmount;
	wire [2:0] bundleOut_0_a_bits_mask_sizeOH = _bundleOut_0_a_bits_mask_sizeOH_T_1[2:0] | 3'h1;
	wire _bundleOut_0_a_bits_mask_T = auto_in_a_bits_size >= 3'h3;
	wire bundleOut_0_a_bits_mask_size = bundleOut_0_a_bits_mask_sizeOH[2];
	wire bundleOut_0_a_bits_mask_bit = auto_in_a_bits_address[2];
	wire bundleOut_0_a_bits_mask_nbit = ~bundleOut_0_a_bits_mask_bit;
	wire bundleOut_0_a_bits_mask_acc = _bundleOut_0_a_bits_mask_T | (bundleOut_0_a_bits_mask_size & bundleOut_0_a_bits_mask_nbit);
	wire bundleOut_0_a_bits_mask_acc_1 = _bundleOut_0_a_bits_mask_T | (bundleOut_0_a_bits_mask_size & bundleOut_0_a_bits_mask_bit);
	wire bundleOut_0_a_bits_mask_size_1 = bundleOut_0_a_bits_mask_sizeOH[1];
	wire bundleOut_0_a_bits_mask_bit_1 = auto_in_a_bits_address[1];
	wire bundleOut_0_a_bits_mask_nbit_1 = ~bundleOut_0_a_bits_mask_bit_1;
	wire bundleOut_0_a_bits_mask_eq_2 = bundleOut_0_a_bits_mask_nbit & bundleOut_0_a_bits_mask_nbit_1;
	wire bundleOut_0_a_bits_mask_acc_2 = bundleOut_0_a_bits_mask_acc | (bundleOut_0_a_bits_mask_size_1 & bundleOut_0_a_bits_mask_eq_2);
	wire bundleOut_0_a_bits_mask_eq_3 = bundleOut_0_a_bits_mask_nbit & bundleOut_0_a_bits_mask_bit_1;
	wire bundleOut_0_a_bits_mask_acc_3 = bundleOut_0_a_bits_mask_acc | (bundleOut_0_a_bits_mask_size_1 & bundleOut_0_a_bits_mask_eq_3);
	wire bundleOut_0_a_bits_mask_eq_4 = bundleOut_0_a_bits_mask_bit & bundleOut_0_a_bits_mask_nbit_1;
	wire bundleOut_0_a_bits_mask_acc_4 = bundleOut_0_a_bits_mask_acc_1 | (bundleOut_0_a_bits_mask_size_1 & bundleOut_0_a_bits_mask_eq_4);
	wire bundleOut_0_a_bits_mask_eq_5 = bundleOut_0_a_bits_mask_bit & bundleOut_0_a_bits_mask_bit_1;
	wire bundleOut_0_a_bits_mask_acc_5 = bundleOut_0_a_bits_mask_acc_1 | (bundleOut_0_a_bits_mask_size_1 & bundleOut_0_a_bits_mask_eq_5);
	wire bundleOut_0_a_bits_mask_size_2 = bundleOut_0_a_bits_mask_sizeOH[0];
	wire bundleOut_0_a_bits_mask_bit_2 = auto_in_a_bits_address[0];
	wire bundleOut_0_a_bits_mask_nbit_2 = ~bundleOut_0_a_bits_mask_bit_2;
	wire bundleOut_0_a_bits_mask_eq_6 = bundleOut_0_a_bits_mask_eq_2 & bundleOut_0_a_bits_mask_nbit_2;
	wire bundleOut_0_a_bits_mask_acc_6 = bundleOut_0_a_bits_mask_acc_2 | (bundleOut_0_a_bits_mask_size_2 & bundleOut_0_a_bits_mask_eq_6);
	wire bundleOut_0_a_bits_mask_eq_7 = bundleOut_0_a_bits_mask_eq_2 & bundleOut_0_a_bits_mask_bit_2;
	wire bundleOut_0_a_bits_mask_acc_7 = bundleOut_0_a_bits_mask_acc_2 | (bundleOut_0_a_bits_mask_size_2 & bundleOut_0_a_bits_mask_eq_7);
	wire bundleOut_0_a_bits_mask_eq_8 = bundleOut_0_a_bits_mask_eq_3 & bundleOut_0_a_bits_mask_nbit_2;
	wire bundleOut_0_a_bits_mask_acc_8 = bundleOut_0_a_bits_mask_acc_3 | (bundleOut_0_a_bits_mask_size_2 & bundleOut_0_a_bits_mask_eq_8);
	wire bundleOut_0_a_bits_mask_eq_9 = bundleOut_0_a_bits_mask_eq_3 & bundleOut_0_a_bits_mask_bit_2;
	wire bundleOut_0_a_bits_mask_acc_9 = bundleOut_0_a_bits_mask_acc_3 | (bundleOut_0_a_bits_mask_size_2 & bundleOut_0_a_bits_mask_eq_9);
	wire bundleOut_0_a_bits_mask_eq_10 = bundleOut_0_a_bits_mask_eq_4 & bundleOut_0_a_bits_mask_nbit_2;
	wire bundleOut_0_a_bits_mask_acc_10 = bundleOut_0_a_bits_mask_acc_4 | (bundleOut_0_a_bits_mask_size_2 & bundleOut_0_a_bits_mask_eq_10);
	wire bundleOut_0_a_bits_mask_eq_11 = bundleOut_0_a_bits_mask_eq_4 & bundleOut_0_a_bits_mask_bit_2;
	wire bundleOut_0_a_bits_mask_acc_11 = bundleOut_0_a_bits_mask_acc_4 | (bundleOut_0_a_bits_mask_size_2 & bundleOut_0_a_bits_mask_eq_11);
	wire bundleOut_0_a_bits_mask_eq_12 = bundleOut_0_a_bits_mask_eq_5 & bundleOut_0_a_bits_mask_nbit_2;
	wire bundleOut_0_a_bits_mask_acc_12 = bundleOut_0_a_bits_mask_acc_5 | (bundleOut_0_a_bits_mask_size_2 & bundleOut_0_a_bits_mask_eq_12);
	wire bundleOut_0_a_bits_mask_eq_13 = bundleOut_0_a_bits_mask_eq_5 & bundleOut_0_a_bits_mask_bit_2;
	wire bundleOut_0_a_bits_mask_acc_13 = bundleOut_0_a_bits_mask_acc_5 | (bundleOut_0_a_bits_mask_size_2 & bundleOut_0_a_bits_mask_eq_13);
	wire [7:0] _bundleOut_0_a_bits_mask_T_1 = {bundleOut_0_a_bits_mask_acc_13, bundleOut_0_a_bits_mask_acc_12, bundleOut_0_a_bits_mask_acc_11, bundleOut_0_a_bits_mask_acc_10, bundleOut_0_a_bits_mask_acc_9, bundleOut_0_a_bits_mask_acc_8, bundleOut_0_a_bits_mask_acc_7, bundleOut_0_a_bits_mask_acc_6};
	reg bundleOut_0_a_bits_mask_rdata_written_once;
	wire bundleOut_0_a_bits_mask_masked_enable_0 = enable_0 | ~bundleOut_0_a_bits_mask_rdata_written_once;
	reg [3:0] bundleOut_0_a_bits_mask_rdata_0;
	wire [3:0] bundleOut_0_a_bits_mask_mdata_0 = (bundleOut_0_a_bits_mask_masked_enable_0 ? auto_in_a_bits_mask : bundleOut_0_a_bits_mask_rdata_0);
	wire _GEN_6 = (_T & _bundleIn_0_a_ready_T) | bundleOut_0_a_bits_mask_rdata_written_once;
	wire [7:0] _bundleOut_0_a_bits_mask_T_5 = {auto_in_a_bits_mask, bundleOut_0_a_bits_mask_mdata_0};
	wire [7:0] _bundleOut_0_a_bits_mask_T_7 = (hasData ? _bundleOut_0_a_bits_mask_T_5 : 8'hff);
	wire [63:0] cated_bits_data = {repeated_repeater_io_deq_bits_data[63:32], auto_out_d_bits_data[31:0]};
	wire [2:0] cated_bits_opcode = repeated_repeater_io_deq_bits_opcode;
	wire repeat_hasData = cated_bits_opcode[0];
	wire [2:0] cated_bits_size = repeated_repeater_io_deq_bits_size;
	wire [9:0] _repeat_limit_T_1 = 10'h007 << cated_bits_size;
	wire [2:0] _repeat_limit_T_3 = ~_repeat_limit_T_1[2:0];
	wire repeat_limit = _repeat_limit_T_3[2];
	reg repeat_count;
	wire repeat_first = ~repeat_count;
	wire repeat_last = (repeat_count == repeat_limit) | ~repeat_hasData;
	wire cated_valid = repeated_repeater_io_deq_valid;
	wire _repeat_T = auto_in_d_ready & cated_valid;
	reg repeat_sel_sel_sources_0;
	reg repeat_sel_sel_sources_1;
	reg repeat_sel_sel_sources_2;
	reg repeat_sel_sel_sources_4;
	wire [2:0] cated_bits_source = repeated_repeater_io_deq_bits_source;
	reg repeat_sel_hold_r;
	wire _GEN_21 = (3'h1 == cated_bits_source ? repeat_sel_sel_sources_1 : repeat_sel_sel_sources_0);
	wire _GEN_22 = (3'h2 == cated_bits_source ? repeat_sel_sel_sources_2 : _GEN_21);
	wire _GEN_23 = (3'h3 == cated_bits_source ? 1'h0 : _GEN_22);
	wire _GEN_24 = (3'h4 == cated_bits_source ? repeat_sel_sel_sources_4 : _GEN_23);
	wire _GEN_25 = (repeat_first ? _GEN_24 : repeat_sel_hold_r);
	wire repeat_sel = _GEN_25 & ~repeat_limit;
	wire repeat_index = repeat_sel | repeat_count;
	wire [31:0] repeat_bundleIn_0_d_bits_data_mux_0 = cated_bits_data[31:0];
	wire [31:0] repeat_bundleIn_0_d_bits_data_mux_1 = cated_bits_data[63:32];
	TLMonitor_10 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Repeater_1 repeated_repeater(
		.clock(repeated_repeater_clock),
		.reset(repeated_repeater_reset),
		.io_repeat(repeated_repeater_io_repeat),
		.io_enq_ready(repeated_repeater_io_enq_ready),
		.io_enq_valid(repeated_repeater_io_enq_valid),
		.io_enq_bits_opcode(repeated_repeater_io_enq_bits_opcode),
		.io_enq_bits_param(repeated_repeater_io_enq_bits_param),
		.io_enq_bits_size(repeated_repeater_io_enq_bits_size),
		.io_enq_bits_source(repeated_repeater_io_enq_bits_source),
		.io_enq_bits_sink(repeated_repeater_io_enq_bits_sink),
		.io_enq_bits_denied(repeated_repeater_io_enq_bits_denied),
		.io_enq_bits_data(repeated_repeater_io_enq_bits_data),
		.io_enq_bits_corrupt(repeated_repeater_io_enq_bits_corrupt),
		.io_deq_ready(repeated_repeater_io_deq_ready),
		.io_deq_valid(repeated_repeater_io_deq_valid),
		.io_deq_bits_opcode(repeated_repeater_io_deq_bits_opcode),
		.io_deq_bits_param(repeated_repeater_io_deq_bits_param),
		.io_deq_bits_size(repeated_repeater_io_deq_bits_size),
		.io_deq_bits_source(repeated_repeater_io_deq_bits_source),
		.io_deq_bits_sink(repeated_repeater_io_deq_bits_sink),
		.io_deq_bits_denied(repeated_repeater_io_deq_bits_denied),
		.io_deq_bits_data(repeated_repeater_io_deq_bits_data),
		.io_deq_bits_corrupt(repeated_repeater_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = auto_out_a_ready | ~last;
	assign auto_in_d_valid = repeated_repeater_io_deq_valid;
	assign auto_in_d_bits_opcode = repeated_repeater_io_deq_bits_opcode;
	assign auto_in_d_bits_param = repeated_repeater_io_deq_bits_param;
	assign auto_in_d_bits_size = repeated_repeater_io_deq_bits_size;
	assign auto_in_d_bits_source = repeated_repeater_io_deq_bits_source;
	assign auto_in_d_bits_sink = repeated_repeater_io_deq_bits_sink;
	assign auto_in_d_bits_denied = repeated_repeater_io_deq_bits_denied;
	assign auto_in_d_bits_data = (repeat_index ? repeat_bundleIn_0_d_bits_data_mux_1 : repeat_bundleIn_0_d_bits_data_mux_0);
	assign auto_in_d_bits_corrupt = repeated_repeater_io_deq_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid & last;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = _bundleOut_0_a_bits_mask_T_1 & _bundleOut_0_a_bits_mask_T_7;
	assign auto_out_a_bits_data = {auto_in_a_bits_data, bundleOut_0_a_bits_data_mdata_0};
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt | corrupt_reg;
	assign auto_out_d_ready = repeated_repeater_io_enq_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_out_a_ready | ~last;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = repeated_repeater_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = repeated_repeater_io_deq_bits_opcode;
	assign monitor_io_in_d_bits_param = repeated_repeater_io_deq_bits_param;
	assign monitor_io_in_d_bits_size = repeated_repeater_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = repeated_repeater_io_deq_bits_source;
	assign monitor_io_in_d_bits_sink = repeated_repeater_io_deq_bits_sink;
	assign monitor_io_in_d_bits_denied = repeated_repeater_io_deq_bits_denied;
	assign monitor_io_in_d_bits_corrupt = repeated_repeater_io_deq_bits_corrupt;
	assign repeated_repeater_clock = clock;
	assign repeated_repeater_reset = reset;
	assign repeated_repeater_io_repeat = ~repeat_last;
	assign repeated_repeater_io_enq_valid = auto_out_d_valid;
	assign repeated_repeater_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign repeated_repeater_io_enq_bits_param = auto_out_d_bits_param;
	assign repeated_repeater_io_enq_bits_size = auto_out_d_bits_size;
	assign repeated_repeater_io_enq_bits_source = auto_out_d_bits_source;
	assign repeated_repeater_io_enq_bits_sink = auto_out_d_bits_sink;
	assign repeated_repeater_io_enq_bits_denied = auto_out_d_bits_denied;
	assign repeated_repeater_io_enq_bits_data = auto_out_d_bits_data;
	assign repeated_repeater_io_enq_bits_corrupt = auto_out_d_bits_corrupt;
	assign repeated_repeater_io_deq_ready = auto_in_d_ready;
	always @(posedge clock) begin
		if (reset)
			count <= 1'h0;
		else if (_T)
			if (last)
				count <= 1'h0;
			else
				count <= count + 1'h1;
		if (reset)
			corrupt_reg <= 1'h0;
		else if (_T)
			if (last)
				corrupt_reg <= 1'h0;
			else
				corrupt_reg <= corrupt_out;
		if (reset)
			bundleOut_0_a_bits_data_rdata_written_once <= 1'h0;
		else
			bundleOut_0_a_bits_data_rdata_written_once <= _GEN_4;
		if (_T & _bundleIn_0_a_ready_T)
			if (bundleOut_0_a_bits_data_masked_enable_0)
				bundleOut_0_a_bits_data_rdata_0 <= auto_in_a_bits_data;
		if (reset)
			bundleOut_0_a_bits_mask_rdata_written_once <= 1'h0;
		else
			bundleOut_0_a_bits_mask_rdata_written_once <= _GEN_6;
		if (_T & _bundleIn_0_a_ready_T)
			if (bundleOut_0_a_bits_mask_masked_enable_0)
				bundleOut_0_a_bits_mask_rdata_0 <= auto_in_a_bits_mask;
		if (reset)
			repeat_count <= 1'h0;
		else if (_repeat_T)
			if (repeat_last)
				repeat_count <= 1'h0;
			else
				repeat_count <= repeat_count + 1'h1;
		if (_T)
			if (3'h0 == auto_in_a_bits_source)
				repeat_sel_sel_sources_0 <= bundleOut_0_a_bits_mask_bit;
		if (_T)
			if (3'h1 == auto_in_a_bits_source)
				repeat_sel_sel_sources_1 <= bundleOut_0_a_bits_mask_bit;
		if (_T)
			if (3'h2 == auto_in_a_bits_source)
				repeat_sel_sel_sources_2 <= bundleOut_0_a_bits_mask_bit;
		if (_T)
			if (3'h4 == auto_in_a_bits_source)
				repeat_sel_sel_sources_4 <= bundleOut_0_a_bits_mask_bit;
		if (repeat_first)
			if (3'h4 == cated_bits_source)
				repeat_sel_hold_r <= repeat_sel_sel_sources_4;
			else if (3'h3 == cated_bits_source)
				repeat_sel_hold_r <= 1'h0;
			else if (3'h2 == cated_bits_source)
				repeat_sel_hold_r <= repeat_sel_sel_sources_2;
			else
				repeat_sel_hold_r <= _GEN_21;
	end
endmodule
module TLInterconnectCoupler_6 (
	clock,
	reset,
	auto_tlserial_manager_crossing_out_a_ready,
	auto_tlserial_manager_crossing_out_a_valid,
	auto_tlserial_manager_crossing_out_a_bits_opcode,
	auto_tlserial_manager_crossing_out_a_bits_param,
	auto_tlserial_manager_crossing_out_a_bits_size,
	auto_tlserial_manager_crossing_out_a_bits_source,
	auto_tlserial_manager_crossing_out_a_bits_address,
	auto_tlserial_manager_crossing_out_a_bits_mask,
	auto_tlserial_manager_crossing_out_a_bits_data,
	auto_tlserial_manager_crossing_out_a_bits_corrupt,
	auto_tlserial_manager_crossing_out_d_ready,
	auto_tlserial_manager_crossing_out_d_valid,
	auto_tlserial_manager_crossing_out_d_bits_opcode,
	auto_tlserial_manager_crossing_out_d_bits_param,
	auto_tlserial_manager_crossing_out_d_bits_size,
	auto_tlserial_manager_crossing_out_d_bits_source,
	auto_tlserial_manager_crossing_out_d_bits_sink,
	auto_tlserial_manager_crossing_out_d_bits_denied,
	auto_tlserial_manager_crossing_out_d_bits_data,
	auto_tlserial_manager_crossing_out_d_bits_corrupt,
	auto_tl_in_a_ready,
	auto_tl_in_a_valid,
	auto_tl_in_a_bits_opcode,
	auto_tl_in_a_bits_param,
	auto_tl_in_a_bits_size,
	auto_tl_in_a_bits_source,
	auto_tl_in_a_bits_address,
	auto_tl_in_a_bits_mask,
	auto_tl_in_a_bits_data,
	auto_tl_in_a_bits_corrupt,
	auto_tl_in_d_ready,
	auto_tl_in_d_valid,
	auto_tl_in_d_bits_opcode,
	auto_tl_in_d_bits_param,
	auto_tl_in_d_bits_size,
	auto_tl_in_d_bits_source,
	auto_tl_in_d_bits_sink,
	auto_tl_in_d_bits_denied,
	auto_tl_in_d_bits_data,
	auto_tl_in_d_bits_corrupt
);
	input clock;
	input reset;
	input auto_tlserial_manager_crossing_out_a_ready;
	output wire auto_tlserial_manager_crossing_out_a_valid;
	output wire [2:0] auto_tlserial_manager_crossing_out_a_bits_opcode;
	output wire [2:0] auto_tlserial_manager_crossing_out_a_bits_param;
	output wire [2:0] auto_tlserial_manager_crossing_out_a_bits_size;
	output wire [2:0] auto_tlserial_manager_crossing_out_a_bits_source;
	output wire [28:0] auto_tlserial_manager_crossing_out_a_bits_address;
	output wire [7:0] auto_tlserial_manager_crossing_out_a_bits_mask;
	output wire [63:0] auto_tlserial_manager_crossing_out_a_bits_data;
	output wire auto_tlserial_manager_crossing_out_a_bits_corrupt;
	output wire auto_tlserial_manager_crossing_out_d_ready;
	input auto_tlserial_manager_crossing_out_d_valid;
	input [2:0] auto_tlserial_manager_crossing_out_d_bits_opcode;
	input [1:0] auto_tlserial_manager_crossing_out_d_bits_param;
	input [2:0] auto_tlserial_manager_crossing_out_d_bits_size;
	input [2:0] auto_tlserial_manager_crossing_out_d_bits_source;
	input auto_tlserial_manager_crossing_out_d_bits_sink;
	input auto_tlserial_manager_crossing_out_d_bits_denied;
	input [63:0] auto_tlserial_manager_crossing_out_d_bits_data;
	input auto_tlserial_manager_crossing_out_d_bits_corrupt;
	output wire auto_tl_in_a_ready;
	input auto_tl_in_a_valid;
	input [2:0] auto_tl_in_a_bits_opcode;
	input [2:0] auto_tl_in_a_bits_param;
	input [2:0] auto_tl_in_a_bits_size;
	input [2:0] auto_tl_in_a_bits_source;
	input [28:0] auto_tl_in_a_bits_address;
	input [3:0] auto_tl_in_a_bits_mask;
	input [31:0] auto_tl_in_a_bits_data;
	input auto_tl_in_a_bits_corrupt;
	input auto_tl_in_d_ready;
	output wire auto_tl_in_d_valid;
	output wire [2:0] auto_tl_in_d_bits_opcode;
	output wire [1:0] auto_tl_in_d_bits_param;
	output wire [2:0] auto_tl_in_d_bits_size;
	output wire [2:0] auto_tl_in_d_bits_source;
	output wire auto_tl_in_d_bits_sink;
	output wire auto_tl_in_d_bits_denied;
	output wire [31:0] auto_tl_in_d_bits_data;
	output wire auto_tl_in_d_bits_corrupt;
	wire shrinker_auto_in_a_ready;
	wire shrinker_auto_in_a_valid;
	wire [2:0] shrinker_auto_in_a_bits_opcode;
	wire [2:0] shrinker_auto_in_a_bits_param;
	wire [2:0] shrinker_auto_in_a_bits_size;
	wire [2:0] shrinker_auto_in_a_bits_source;
	wire [28:0] shrinker_auto_in_a_bits_address;
	wire [7:0] shrinker_auto_in_a_bits_mask;
	wire [63:0] shrinker_auto_in_a_bits_data;
	wire shrinker_auto_in_a_bits_corrupt;
	wire shrinker_auto_in_d_ready;
	wire shrinker_auto_in_d_valid;
	wire [2:0] shrinker_auto_in_d_bits_opcode;
	wire [1:0] shrinker_auto_in_d_bits_param;
	wire [2:0] shrinker_auto_in_d_bits_size;
	wire [2:0] shrinker_auto_in_d_bits_source;
	wire shrinker_auto_in_d_bits_sink;
	wire shrinker_auto_in_d_bits_denied;
	wire [63:0] shrinker_auto_in_d_bits_data;
	wire shrinker_auto_in_d_bits_corrupt;
	wire shrinker_auto_out_a_ready;
	wire shrinker_auto_out_a_valid;
	wire [2:0] shrinker_auto_out_a_bits_opcode;
	wire [2:0] shrinker_auto_out_a_bits_param;
	wire [2:0] shrinker_auto_out_a_bits_size;
	wire [2:0] shrinker_auto_out_a_bits_source;
	wire [28:0] shrinker_auto_out_a_bits_address;
	wire [7:0] shrinker_auto_out_a_bits_mask;
	wire [63:0] shrinker_auto_out_a_bits_data;
	wire shrinker_auto_out_a_bits_corrupt;
	wire shrinker_auto_out_d_ready;
	wire shrinker_auto_out_d_valid;
	wire [2:0] shrinker_auto_out_d_bits_opcode;
	wire [1:0] shrinker_auto_out_d_bits_param;
	wire [2:0] shrinker_auto_out_d_bits_size;
	wire [2:0] shrinker_auto_out_d_bits_source;
	wire shrinker_auto_out_d_bits_sink;
	wire shrinker_auto_out_d_bits_denied;
	wire [63:0] shrinker_auto_out_d_bits_data;
	wire shrinker_auto_out_d_bits_corrupt;
	wire widget_clock;
	wire widget_reset;
	wire widget_auto_in_a_ready;
	wire widget_auto_in_a_valid;
	wire [2:0] widget_auto_in_a_bits_opcode;
	wire [2:0] widget_auto_in_a_bits_param;
	wire [2:0] widget_auto_in_a_bits_size;
	wire [2:0] widget_auto_in_a_bits_source;
	wire [28:0] widget_auto_in_a_bits_address;
	wire [3:0] widget_auto_in_a_bits_mask;
	wire [31:0] widget_auto_in_a_bits_data;
	wire widget_auto_in_a_bits_corrupt;
	wire widget_auto_in_d_ready;
	wire widget_auto_in_d_valid;
	wire [2:0] widget_auto_in_d_bits_opcode;
	wire [1:0] widget_auto_in_d_bits_param;
	wire [2:0] widget_auto_in_d_bits_size;
	wire [2:0] widget_auto_in_d_bits_source;
	wire widget_auto_in_d_bits_sink;
	wire widget_auto_in_d_bits_denied;
	wire [31:0] widget_auto_in_d_bits_data;
	wire widget_auto_in_d_bits_corrupt;
	wire widget_auto_out_a_ready;
	wire widget_auto_out_a_valid;
	wire [2:0] widget_auto_out_a_bits_opcode;
	wire [2:0] widget_auto_out_a_bits_param;
	wire [2:0] widget_auto_out_a_bits_size;
	wire [2:0] widget_auto_out_a_bits_source;
	wire [28:0] widget_auto_out_a_bits_address;
	wire [7:0] widget_auto_out_a_bits_mask;
	wire [63:0] widget_auto_out_a_bits_data;
	wire widget_auto_out_a_bits_corrupt;
	wire widget_auto_out_d_ready;
	wire widget_auto_out_d_valid;
	wire [2:0] widget_auto_out_d_bits_opcode;
	wire [1:0] widget_auto_out_d_bits_param;
	wire [2:0] widget_auto_out_d_bits_size;
	wire [2:0] widget_auto_out_d_bits_source;
	wire widget_auto_out_d_bits_sink;
	wire widget_auto_out_d_bits_denied;
	wire [63:0] widget_auto_out_d_bits_data;
	wire widget_auto_out_d_bits_corrupt;
	TLSourceShrinker_1 shrinker(
		.auto_in_a_ready(shrinker_auto_in_a_ready),
		.auto_in_a_valid(shrinker_auto_in_a_valid),
		.auto_in_a_bits_opcode(shrinker_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(shrinker_auto_in_a_bits_param),
		.auto_in_a_bits_size(shrinker_auto_in_a_bits_size),
		.auto_in_a_bits_source(shrinker_auto_in_a_bits_source),
		.auto_in_a_bits_address(shrinker_auto_in_a_bits_address),
		.auto_in_a_bits_mask(shrinker_auto_in_a_bits_mask),
		.auto_in_a_bits_data(shrinker_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(shrinker_auto_in_a_bits_corrupt),
		.auto_in_d_ready(shrinker_auto_in_d_ready),
		.auto_in_d_valid(shrinker_auto_in_d_valid),
		.auto_in_d_bits_opcode(shrinker_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(shrinker_auto_in_d_bits_param),
		.auto_in_d_bits_size(shrinker_auto_in_d_bits_size),
		.auto_in_d_bits_source(shrinker_auto_in_d_bits_source),
		.auto_in_d_bits_sink(shrinker_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(shrinker_auto_in_d_bits_denied),
		.auto_in_d_bits_data(shrinker_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(shrinker_auto_in_d_bits_corrupt),
		.auto_out_a_ready(shrinker_auto_out_a_ready),
		.auto_out_a_valid(shrinker_auto_out_a_valid),
		.auto_out_a_bits_opcode(shrinker_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(shrinker_auto_out_a_bits_param),
		.auto_out_a_bits_size(shrinker_auto_out_a_bits_size),
		.auto_out_a_bits_source(shrinker_auto_out_a_bits_source),
		.auto_out_a_bits_address(shrinker_auto_out_a_bits_address),
		.auto_out_a_bits_mask(shrinker_auto_out_a_bits_mask),
		.auto_out_a_bits_data(shrinker_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(shrinker_auto_out_a_bits_corrupt),
		.auto_out_d_ready(shrinker_auto_out_d_ready),
		.auto_out_d_valid(shrinker_auto_out_d_valid),
		.auto_out_d_bits_opcode(shrinker_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(shrinker_auto_out_d_bits_param),
		.auto_out_d_bits_size(shrinker_auto_out_d_bits_size),
		.auto_out_d_bits_source(shrinker_auto_out_d_bits_source),
		.auto_out_d_bits_sink(shrinker_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(shrinker_auto_out_d_bits_denied),
		.auto_out_d_bits_data(shrinker_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(shrinker_auto_out_d_bits_corrupt)
	);
	TLWidthWidget_4 widget(
		.clock(widget_clock),
		.reset(widget_reset),
		.auto_in_a_ready(widget_auto_in_a_ready),
		.auto_in_a_valid(widget_auto_in_a_valid),
		.auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(widget_auto_in_a_bits_param),
		.auto_in_a_bits_size(widget_auto_in_a_bits_size),
		.auto_in_a_bits_source(widget_auto_in_a_bits_source),
		.auto_in_a_bits_address(widget_auto_in_a_bits_address),
		.auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
		.auto_in_a_bits_data(widget_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(widget_auto_in_a_bits_corrupt),
		.auto_in_d_ready(widget_auto_in_d_ready),
		.auto_in_d_valid(widget_auto_in_d_valid),
		.auto_in_d_bits_opcode(widget_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(widget_auto_in_d_bits_param),
		.auto_in_d_bits_size(widget_auto_in_d_bits_size),
		.auto_in_d_bits_source(widget_auto_in_d_bits_source),
		.auto_in_d_bits_sink(widget_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(widget_auto_in_d_bits_denied),
		.auto_in_d_bits_data(widget_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(widget_auto_in_d_bits_corrupt),
		.auto_out_a_ready(widget_auto_out_a_ready),
		.auto_out_a_valid(widget_auto_out_a_valid),
		.auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(widget_auto_out_a_bits_param),
		.auto_out_a_bits_size(widget_auto_out_a_bits_size),
		.auto_out_a_bits_source(widget_auto_out_a_bits_source),
		.auto_out_a_bits_address(widget_auto_out_a_bits_address),
		.auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
		.auto_out_a_bits_data(widget_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(widget_auto_out_a_bits_corrupt),
		.auto_out_d_ready(widget_auto_out_d_ready),
		.auto_out_d_valid(widget_auto_out_d_valid),
		.auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(widget_auto_out_d_bits_param),
		.auto_out_d_bits_size(widget_auto_out_d_bits_size),
		.auto_out_d_bits_source(widget_auto_out_d_bits_source),
		.auto_out_d_bits_sink(widget_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(widget_auto_out_d_bits_denied),
		.auto_out_d_bits_data(widget_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(widget_auto_out_d_bits_corrupt)
	);
	assign auto_tlserial_manager_crossing_out_a_valid = shrinker_auto_out_a_valid;
	assign auto_tlserial_manager_crossing_out_a_bits_opcode = shrinker_auto_out_a_bits_opcode;
	assign auto_tlserial_manager_crossing_out_a_bits_param = shrinker_auto_out_a_bits_param;
	assign auto_tlserial_manager_crossing_out_a_bits_size = shrinker_auto_out_a_bits_size;
	assign auto_tlserial_manager_crossing_out_a_bits_source = shrinker_auto_out_a_bits_source;
	assign auto_tlserial_manager_crossing_out_a_bits_address = shrinker_auto_out_a_bits_address;
	assign auto_tlserial_manager_crossing_out_a_bits_mask = shrinker_auto_out_a_bits_mask;
	assign auto_tlserial_manager_crossing_out_a_bits_data = shrinker_auto_out_a_bits_data;
	assign auto_tlserial_manager_crossing_out_a_bits_corrupt = shrinker_auto_out_a_bits_corrupt;
	assign auto_tlserial_manager_crossing_out_d_ready = shrinker_auto_out_d_ready;
	assign auto_tl_in_a_ready = widget_auto_in_a_ready;
	assign auto_tl_in_d_valid = widget_auto_in_d_valid;
	assign auto_tl_in_d_bits_opcode = widget_auto_in_d_bits_opcode;
	assign auto_tl_in_d_bits_param = widget_auto_in_d_bits_param;
	assign auto_tl_in_d_bits_size = widget_auto_in_d_bits_size;
	assign auto_tl_in_d_bits_source = widget_auto_in_d_bits_source;
	assign auto_tl_in_d_bits_sink = widget_auto_in_d_bits_sink;
	assign auto_tl_in_d_bits_denied = widget_auto_in_d_bits_denied;
	assign auto_tl_in_d_bits_data = widget_auto_in_d_bits_data;
	assign auto_tl_in_d_bits_corrupt = widget_auto_in_d_bits_corrupt;
	assign shrinker_auto_in_a_valid = widget_auto_out_a_valid;
	assign shrinker_auto_in_a_bits_opcode = widget_auto_out_a_bits_opcode;
	assign shrinker_auto_in_a_bits_param = widget_auto_out_a_bits_param;
	assign shrinker_auto_in_a_bits_size = widget_auto_out_a_bits_size;
	assign shrinker_auto_in_a_bits_source = widget_auto_out_a_bits_source;
	assign shrinker_auto_in_a_bits_address = widget_auto_out_a_bits_address;
	assign shrinker_auto_in_a_bits_mask = widget_auto_out_a_bits_mask;
	assign shrinker_auto_in_a_bits_data = widget_auto_out_a_bits_data;
	assign shrinker_auto_in_a_bits_corrupt = widget_auto_out_a_bits_corrupt;
	assign shrinker_auto_in_d_ready = widget_auto_out_d_ready;
	assign shrinker_auto_out_a_ready = auto_tlserial_manager_crossing_out_a_ready;
	assign shrinker_auto_out_d_valid = auto_tlserial_manager_crossing_out_d_valid;
	assign shrinker_auto_out_d_bits_opcode = auto_tlserial_manager_crossing_out_d_bits_opcode;
	assign shrinker_auto_out_d_bits_param = auto_tlserial_manager_crossing_out_d_bits_param;
	assign shrinker_auto_out_d_bits_size = auto_tlserial_manager_crossing_out_d_bits_size;
	assign shrinker_auto_out_d_bits_source = auto_tlserial_manager_crossing_out_d_bits_source;
	assign shrinker_auto_out_d_bits_sink = auto_tlserial_manager_crossing_out_d_bits_sink;
	assign shrinker_auto_out_d_bits_denied = auto_tlserial_manager_crossing_out_d_bits_denied;
	assign shrinker_auto_out_d_bits_data = auto_tlserial_manager_crossing_out_d_bits_data;
	assign shrinker_auto_out_d_bits_corrupt = auto_tlserial_manager_crossing_out_d_bits_corrupt;
	assign widget_clock = clock;
	assign widget_reset = reset;
	assign widget_auto_in_a_valid = auto_tl_in_a_valid;
	assign widget_auto_in_a_bits_opcode = auto_tl_in_a_bits_opcode;
	assign widget_auto_in_a_bits_param = auto_tl_in_a_bits_param;
	assign widget_auto_in_a_bits_size = auto_tl_in_a_bits_size;
	assign widget_auto_in_a_bits_source = auto_tl_in_a_bits_source;
	assign widget_auto_in_a_bits_address = auto_tl_in_a_bits_address;
	assign widget_auto_in_a_bits_mask = auto_tl_in_a_bits_mask;
	assign widget_auto_in_a_bits_data = auto_tl_in_a_bits_data;
	assign widget_auto_in_a_bits_corrupt = auto_tl_in_a_bits_corrupt;
	assign widget_auto_in_d_ready = auto_tl_in_d_ready;
	assign widget_auto_out_a_ready = shrinker_auto_in_a_ready;
	assign widget_auto_out_d_valid = shrinker_auto_in_d_valid;
	assign widget_auto_out_d_bits_opcode = shrinker_auto_in_d_bits_opcode;
	assign widget_auto_out_d_bits_param = shrinker_auto_in_d_bits_param;
	assign widget_auto_out_d_bits_size = shrinker_auto_in_d_bits_size;
	assign widget_auto_out_d_bits_source = shrinker_auto_in_d_bits_source;
	assign widget_auto_out_d_bits_sink = shrinker_auto_in_d_bits_sink;
	assign widget_auto_out_d_bits_denied = shrinker_auto_in_d_bits_denied;
	assign widget_auto_out_d_bits_data = shrinker_auto_in_d_bits_data;
	assign widget_auto_out_d_bits_corrupt = shrinker_auto_in_d_bits_corrupt;
endmodule
module TLMonitor_11 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [30:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [30:0] _GEN_71 = {25'd0, is_aligned_mask};
	wire [30:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 31'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [30:0] _T_56 = io_in_a_bits_address ^ 31'h54000000;
	wire [31:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [31:0] _T_59 = $signed(_T_57) & -32'sh00001000;
	wire _T_60 = $signed(_T_59) == 32'sh00000000;
	wire _T_92 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_96 = ~io_in_a_bits_mask;
	wire _T_97 = _T_96 == 4'h0;
	wire _T_101 = ~io_in_a_bits_corrupt;
	wire _T_105 = io_in_a_bits_opcode == 3'h7;
	wire _T_159 = io_in_a_bits_param != 3'h0;
	wire _T_172 = io_in_a_bits_opcode == 3'h4;
	wire _T_189 = io_in_a_bits_size <= 3'h6;
	wire _T_197 = _T_189 & _T_60;
	wire _T_208 = io_in_a_bits_param == 3'h0;
	wire _T_212 = io_in_a_bits_mask == mask;
	wire _T_220 = io_in_a_bits_opcode == 3'h0;
	wire _T_244 = source_ok & _T_197;
	wire _T_262 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_300 = ~mask;
	wire [3:0] _T_301 = io_in_a_bits_mask & _T_300;
	wire _T_302 = _T_301 == 4'h0;
	wire _T_306 = io_in_a_bits_opcode == 3'h2;
	wire _T_337 = io_in_a_bits_param <= 3'h4;
	wire _T_345 = io_in_a_bits_opcode == 3'h3;
	wire _T_376 = io_in_a_bits_param <= 3'h3;
	wire _T_384 = io_in_a_bits_opcode == 3'h5;
	wire _T_415 = io_in_a_bits_param <= 3'h1;
	wire _T_427 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_431 = io_in_d_bits_opcode == 3'h6;
	wire _T_435 = io_in_d_bits_size >= 3'h2;
	wire _T_451 = io_in_d_bits_opcode == 3'h4;
	wire _T_479 = io_in_d_bits_opcode == 3'h5;
	wire _T_508 = io_in_d_bits_opcode == 3'h0;
	wire _T_525 = io_in_d_bits_opcode == 3'h1;
	wire _T_543 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [30:0] address;
	wire _T_573 = io_in_a_valid & ~a_first;
	wire _T_574 = io_in_a_bits_opcode == opcode;
	wire _T_578 = io_in_a_bits_param == param;
	wire _T_582 = io_in_a_bits_size == size;
	wire _T_586 = io_in_a_bits_source == source;
	wire _T_590 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	wire _T_597 = io_in_d_valid & ~d_first;
	wire _T_598 = io_in_d_bits_opcode == opcode_1;
	wire _T_606 = io_in_d_bits_size == size_1;
	wire _T_610 = io_in_d_bits_source == source_1;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_624 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire _T_627 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_629 = inflight >> io_in_a_bits_source;
	wire _T_631 = ~_T_629[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_635 = io_in_d_valid & d_first_1;
	wire _T_637 = ~_T_431;
	wire _T_638 = (io_in_d_valid & d_first_1) & ~_T_431;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_637 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_637 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_624 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_648 = inflight >> io_in_d_bits_source;
	wire _T_650 = _T_648[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_655 = io_in_d_bits_opcode == _GEN_40;
	wire _T_656 = (io_in_d_bits_opcode == _GEN_32) | _T_655;
	wire _T_660 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_667 = io_in_d_bits_opcode == _GEN_56;
	wire _T_668 = (io_in_d_bits_opcode == _GEN_48) | _T_667;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_672 = _GEN_82 == a_size_lookup;
	wire _T_682 = (((_T_635 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_637;
	wire _T_684 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_693 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_719 = (io_in_d_valid & d_first_2) & _T_431;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_431 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_431 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_727 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_737 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_757 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Repeater_2 (
	clock,
	reset,
	io_repeat,
	io_full,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	input io_repeat;
	output wire io_full;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [30:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [30:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire io_deq_bits_corrupt;
	reg full;
	reg [2:0] saved_opcode;
	reg [2:0] saved_param;
	reg [2:0] saved_size;
	reg [2:0] saved_source;
	reg [30:0] saved_address;
	reg [3:0] saved_mask;
	reg saved_corrupt;
	wire _T = io_enq_ready & io_enq_valid;
	wire _GEN_0 = (_T & io_repeat) | full;
	wire _T_2 = io_deq_ready & io_deq_valid;
	assign io_full = full;
	assign io_enq_ready = io_deq_ready & ~full;
	assign io_deq_valid = io_enq_valid | full;
	assign io_deq_bits_opcode = (full ? saved_opcode : io_enq_bits_opcode);
	assign io_deq_bits_param = (full ? saved_param : io_enq_bits_param);
	assign io_deq_bits_size = (full ? saved_size : io_enq_bits_size);
	assign io_deq_bits_source = (full ? saved_source : io_enq_bits_source);
	assign io_deq_bits_address = (full ? saved_address : io_enq_bits_address);
	assign io_deq_bits_mask = (full ? saved_mask : io_enq_bits_mask);
	assign io_deq_bits_corrupt = (full ? saved_corrupt : io_enq_bits_corrupt);
	always @(posedge clock) begin
		if (reset)
			full <= 1'h0;
		else if (_T_2 & ~io_repeat)
			full <= 1'h0;
		else
			full <= _GEN_0;
		if (_T & io_repeat)
			saved_opcode <= io_enq_bits_opcode;
		if (_T & io_repeat)
			saved_param <= io_enq_bits_param;
		if (_T & io_repeat)
			saved_size <= io_enq_bits_size;
		if (_T & io_repeat)
			saved_source <= io_enq_bits_source;
		if (_T & io_repeat)
			saved_address <= io_enq_bits_address;
		if (_T & io_repeat)
			saved_mask <= io_enq_bits_mask;
		if (_T & io_repeat)
			saved_corrupt <= io_enq_bits_corrupt;
	end
endmodule
module TLFragmenter_1 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [30:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire [7:0] auto_out_a_bits_source;
	output wire [30:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_size;
	input [7:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [30:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire repeater_clock;
	wire repeater_reset;
	wire repeater_io_repeat;
	wire repeater_io_full;
	wire repeater_io_enq_ready;
	wire repeater_io_enq_valid;
	wire [2:0] repeater_io_enq_bits_opcode;
	wire [2:0] repeater_io_enq_bits_param;
	wire [2:0] repeater_io_enq_bits_size;
	wire [2:0] repeater_io_enq_bits_source;
	wire [30:0] repeater_io_enq_bits_address;
	wire [3:0] repeater_io_enq_bits_mask;
	wire repeater_io_enq_bits_corrupt;
	wire repeater_io_deq_ready;
	wire repeater_io_deq_valid;
	wire [2:0] repeater_io_deq_bits_opcode;
	wire [2:0] repeater_io_deq_bits_param;
	wire [2:0] repeater_io_deq_bits_size;
	wire [2:0] repeater_io_deq_bits_source;
	wire [30:0] repeater_io_deq_bits_address;
	wire [3:0] repeater_io_deq_bits_mask;
	wire repeater_io_deq_bits_corrupt;
	reg [3:0] acknum;
	reg [2:0] dOrig;
	reg dToggle;
	wire [3:0] dFragnum = auto_out_d_bits_source[3:0];
	wire dFirst = acknum == 4'h0;
	wire dLast = dFragnum == 4'h0;
	wire [3:0] _dsizeOH_T = 4'h1 << auto_out_d_bits_size;
	wire [2:0] dsizeOH = _dsizeOH_T[2:0];
	wire [4:0] _dsizeOH1_T_1 = 5'h03 << auto_out_d_bits_size;
	wire [1:0] dsizeOH1 = ~_dsizeOH1_T_1[1:0];
	wire dHasData = auto_out_d_bits_opcode[0];
	wire _T_5 = ~reset;
	wire ack_decrement = dHasData | dsizeOH[2];
	wire [5:0] _dFirst_size_T = {dFragnum, 2'h0};
	wire [5:0] _GEN_7 = {4'd0, dsizeOH1};
	wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7;
	wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0};
	wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h01;
	wire [6:0] _dFirst_size_T_4 = {1'h0, _dFirst_size_T_1};
	wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4;
	wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5;
	wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4];
	wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0];
	wire _dFirst_size_T_7 = |dFirst_size_hi;
	wire [3:0] _GEN_8 = {1'd0, dFirst_size_hi};
	wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo;
	wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2];
	wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0];
	wire _dFirst_size_T_9 = |dFirst_size_hi_1;
	wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1;
	wire [2:0] dFirst_size = {_dFirst_size_T_7, _dFirst_size_T_9, _dFirst_size_T_10[1]};
	wire drop = ~dHasData & ~dLast;
	wire bundleOut_0_d_ready = auto_in_d_ready | drop;
	wire _T_7 = bundleOut_0_d_ready & auto_out_d_valid;
	wire [3:0] _GEN_9 = {3'd0, ack_decrement};
	wire [3:0] _acknum_T_1 = acknum - _GEN_9;
	wire [2:0] aFrag = (repeater_io_deq_bits_size > 3'h2 ? 3'h2 : repeater_io_deq_bits_size);
	wire [12:0] _aOrigOH1_T_1 = 13'h003f << repeater_io_deq_bits_size;
	wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0];
	wire [8:0] _aFragOH1_T_1 = 9'h003 << aFrag;
	wire [1:0] aFragOH1 = ~_aFragOH1_T_1[1:0];
	wire aHasData = ~repeater_io_deq_bits_opcode[2];
	reg [3:0] gennum;
	wire aFirst = gennum == 4'h0;
	wire [3:0] _old_gennum1_T_2 = gennum - 4'h1;
	wire [3:0] old_gennum1 = (aFirst ? aOrigOH1[5:2] : _old_gennum1_T_2);
	wire [3:0] _new_gennum_T = ~old_gennum1;
	wire [3:0] new_gennum = ~_new_gennum_T;
	reg aToggle_r;
	wire _GEN_5 = (aFirst ? dToggle : aToggle_r);
	wire aToggle = ~_GEN_5;
	wire bundleOut_0_a_valid = repeater_io_deq_valid;
	wire _T_8 = auto_out_a_ready & bundleOut_0_a_valid;
	wire _repeater_io_repeat_T = ~aHasData;
	wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 2'h0};
	wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1;
	wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1;
	wire [5:0] _GEN_10 = {4'd0, aFragOH1};
	wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10;
	wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h03;
	wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4;
	wire [30:0] _GEN_11 = {25'd0, _bundleOut_0_a_bits_address_T_5};
	wire [3:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source, aToggle};
	wire _T_9 = ~repeater_io_full;
	TLMonitor_11 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	Repeater_2 repeater(
		.clock(repeater_clock),
		.reset(repeater_reset),
		.io_repeat(repeater_io_repeat),
		.io_full(repeater_io_full),
		.io_enq_ready(repeater_io_enq_ready),
		.io_enq_valid(repeater_io_enq_valid),
		.io_enq_bits_opcode(repeater_io_enq_bits_opcode),
		.io_enq_bits_param(repeater_io_enq_bits_param),
		.io_enq_bits_size(repeater_io_enq_bits_size),
		.io_enq_bits_source(repeater_io_enq_bits_source),
		.io_enq_bits_address(repeater_io_enq_bits_address),
		.io_enq_bits_mask(repeater_io_enq_bits_mask),
		.io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
		.io_deq_ready(repeater_io_deq_ready),
		.io_deq_valid(repeater_io_deq_valid),
		.io_deq_bits_opcode(repeater_io_deq_bits_opcode),
		.io_deq_bits_param(repeater_io_deq_bits_param),
		.io_deq_bits_size(repeater_io_deq_bits_size),
		.io_deq_bits_source(repeater_io_deq_bits_source),
		.io_deq_bits_address(repeater_io_deq_bits_address),
		.io_deq_bits_mask(repeater_io_deq_bits_mask),
		.io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = repeater_io_enq_ready;
	assign auto_in_d_valid = auto_out_d_valid & ~drop;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign auto_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_out_a_valid = repeater_io_deq_valid;
	assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode;
	assign auto_out_a_bits_param = repeater_io_deq_bits_param;
	assign auto_out_a_bits_size = aFrag[1:0];
	assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi, new_gennum};
	assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11;
	assign auto_out_a_bits_mask = (repeater_io_full ? 4'hf : auto_in_a_bits_mask);
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready | drop;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = repeater_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid & ~drop;
	assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_io_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign repeater_clock = clock;
	assign repeater_reset = reset;
	assign repeater_io_repeat = ~aHasData & (new_gennum != 4'h0);
	assign repeater_io_enq_valid = auto_in_a_valid;
	assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign repeater_io_enq_bits_param = auto_in_a_bits_param;
	assign repeater_io_enq_bits_size = auto_in_a_bits_size;
	assign repeater_io_enq_bits_source = auto_in_a_bits_source;
	assign repeater_io_enq_bits_address = auto_in_a_bits_address;
	assign repeater_io_enq_bits_mask = auto_in_a_bits_mask;
	assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign repeater_io_deq_ready = auto_out_a_ready;
	always @(posedge clock) begin
		if (reset)
			acknum <= 4'h0;
		else if (_T_7)
			if (dFirst)
				acknum <= dFragnum;
			else
				acknum <= _acknum_T_1;
		if (_T_7)
			if (dFirst)
				dOrig <= dFirst_size;
		if (reset)
			dToggle <= 1'h0;
		else if (_T_7)
			if (dFirst)
				dToggle <= auto_out_d_bits_source[4];
		if (reset)
			gennum <= 4'h0;
		else if (_T_8)
			gennum <= new_gennum;
		if (aFirst)
			aToggle_r <= dToggle;
	end
endmodule
module TLInterconnectCoupler_7 (
	clock,
	reset,
	auto_control_xing_out_a_ready,
	auto_control_xing_out_a_valid,
	auto_control_xing_out_a_bits_opcode,
	auto_control_xing_out_a_bits_param,
	auto_control_xing_out_a_bits_size,
	auto_control_xing_out_a_bits_source,
	auto_control_xing_out_a_bits_address,
	auto_control_xing_out_a_bits_mask,
	auto_control_xing_out_a_bits_data,
	auto_control_xing_out_a_bits_corrupt,
	auto_control_xing_out_d_ready,
	auto_control_xing_out_d_valid,
	auto_control_xing_out_d_bits_opcode,
	auto_control_xing_out_d_bits_size,
	auto_control_xing_out_d_bits_source,
	auto_control_xing_out_d_bits_data,
	auto_tl_in_a_ready,
	auto_tl_in_a_valid,
	auto_tl_in_a_bits_opcode,
	auto_tl_in_a_bits_param,
	auto_tl_in_a_bits_size,
	auto_tl_in_a_bits_source,
	auto_tl_in_a_bits_address,
	auto_tl_in_a_bits_mask,
	auto_tl_in_a_bits_data,
	auto_tl_in_a_bits_corrupt,
	auto_tl_in_d_ready,
	auto_tl_in_d_valid,
	auto_tl_in_d_bits_opcode,
	auto_tl_in_d_bits_size,
	auto_tl_in_d_bits_source,
	auto_tl_in_d_bits_data
);
	input clock;
	input reset;
	input auto_control_xing_out_a_ready;
	output wire auto_control_xing_out_a_valid;
	output wire [2:0] auto_control_xing_out_a_bits_opcode;
	output wire [2:0] auto_control_xing_out_a_bits_param;
	output wire [1:0] auto_control_xing_out_a_bits_size;
	output wire [7:0] auto_control_xing_out_a_bits_source;
	output wire [30:0] auto_control_xing_out_a_bits_address;
	output wire [3:0] auto_control_xing_out_a_bits_mask;
	output wire [31:0] auto_control_xing_out_a_bits_data;
	output wire auto_control_xing_out_a_bits_corrupt;
	output wire auto_control_xing_out_d_ready;
	input auto_control_xing_out_d_valid;
	input [2:0] auto_control_xing_out_d_bits_opcode;
	input [1:0] auto_control_xing_out_d_bits_size;
	input [7:0] auto_control_xing_out_d_bits_source;
	input [31:0] auto_control_xing_out_d_bits_data;
	output wire auto_tl_in_a_ready;
	input auto_tl_in_a_valid;
	input [2:0] auto_tl_in_a_bits_opcode;
	input [2:0] auto_tl_in_a_bits_param;
	input [2:0] auto_tl_in_a_bits_size;
	input [2:0] auto_tl_in_a_bits_source;
	input [30:0] auto_tl_in_a_bits_address;
	input [3:0] auto_tl_in_a_bits_mask;
	input [31:0] auto_tl_in_a_bits_data;
	input auto_tl_in_a_bits_corrupt;
	input auto_tl_in_d_ready;
	output wire auto_tl_in_d_valid;
	output wire [2:0] auto_tl_in_d_bits_opcode;
	output wire [2:0] auto_tl_in_d_bits_size;
	output wire [2:0] auto_tl_in_d_bits_source;
	output wire [31:0] auto_tl_in_d_bits_data;
	wire fragmenter_clock;
	wire fragmenter_reset;
	wire fragmenter_auto_in_a_ready;
	wire fragmenter_auto_in_a_valid;
	wire [2:0] fragmenter_auto_in_a_bits_opcode;
	wire [2:0] fragmenter_auto_in_a_bits_param;
	wire [2:0] fragmenter_auto_in_a_bits_size;
	wire [2:0] fragmenter_auto_in_a_bits_source;
	wire [30:0] fragmenter_auto_in_a_bits_address;
	wire [3:0] fragmenter_auto_in_a_bits_mask;
	wire [31:0] fragmenter_auto_in_a_bits_data;
	wire fragmenter_auto_in_a_bits_corrupt;
	wire fragmenter_auto_in_d_ready;
	wire fragmenter_auto_in_d_valid;
	wire [2:0] fragmenter_auto_in_d_bits_opcode;
	wire [2:0] fragmenter_auto_in_d_bits_size;
	wire [2:0] fragmenter_auto_in_d_bits_source;
	wire [31:0] fragmenter_auto_in_d_bits_data;
	wire fragmenter_auto_out_a_ready;
	wire fragmenter_auto_out_a_valid;
	wire [2:0] fragmenter_auto_out_a_bits_opcode;
	wire [2:0] fragmenter_auto_out_a_bits_param;
	wire [1:0] fragmenter_auto_out_a_bits_size;
	wire [7:0] fragmenter_auto_out_a_bits_source;
	wire [30:0] fragmenter_auto_out_a_bits_address;
	wire [3:0] fragmenter_auto_out_a_bits_mask;
	wire [31:0] fragmenter_auto_out_a_bits_data;
	wire fragmenter_auto_out_a_bits_corrupt;
	wire fragmenter_auto_out_d_ready;
	wire fragmenter_auto_out_d_valid;
	wire [2:0] fragmenter_auto_out_d_bits_opcode;
	wire [1:0] fragmenter_auto_out_d_bits_size;
	wire [7:0] fragmenter_auto_out_d_bits_source;
	wire [31:0] fragmenter_auto_out_d_bits_data;
	TLFragmenter_1 fragmenter(
		.clock(fragmenter_clock),
		.reset(fragmenter_reset),
		.auto_in_a_ready(fragmenter_auto_in_a_ready),
		.auto_in_a_valid(fragmenter_auto_in_a_valid),
		.auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
		.auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
		.auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
		.auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
		.auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
		.auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
		.auto_in_d_ready(fragmenter_auto_in_d_ready),
		.auto_in_d_valid(fragmenter_auto_in_d_valid),
		.auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
		.auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
		.auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
		.auto_out_a_ready(fragmenter_auto_out_a_ready),
		.auto_out_a_valid(fragmenter_auto_out_a_valid),
		.auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
		.auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
		.auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
		.auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
		.auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
		.auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
		.auto_out_d_ready(fragmenter_auto_out_d_ready),
		.auto_out_d_valid(fragmenter_auto_out_d_valid),
		.auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
		.auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
		.auto_out_d_bits_data(fragmenter_auto_out_d_bits_data)
	);
	assign auto_control_xing_out_a_valid = fragmenter_auto_out_a_valid;
	assign auto_control_xing_out_a_bits_opcode = fragmenter_auto_out_a_bits_opcode;
	assign auto_control_xing_out_a_bits_param = fragmenter_auto_out_a_bits_param;
	assign auto_control_xing_out_a_bits_size = fragmenter_auto_out_a_bits_size;
	assign auto_control_xing_out_a_bits_source = fragmenter_auto_out_a_bits_source;
	assign auto_control_xing_out_a_bits_address = fragmenter_auto_out_a_bits_address;
	assign auto_control_xing_out_a_bits_mask = fragmenter_auto_out_a_bits_mask;
	assign auto_control_xing_out_a_bits_data = fragmenter_auto_out_a_bits_data;
	assign auto_control_xing_out_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt;
	assign auto_control_xing_out_d_ready = fragmenter_auto_out_d_ready;
	assign auto_tl_in_a_ready = fragmenter_auto_in_a_ready;
	assign auto_tl_in_d_valid = fragmenter_auto_in_d_valid;
	assign auto_tl_in_d_bits_opcode = fragmenter_auto_in_d_bits_opcode;
	assign auto_tl_in_d_bits_size = fragmenter_auto_in_d_bits_size;
	assign auto_tl_in_d_bits_source = fragmenter_auto_in_d_bits_source;
	assign auto_tl_in_d_bits_data = fragmenter_auto_in_d_bits_data;
	assign fragmenter_clock = clock;
	assign fragmenter_reset = reset;
	assign fragmenter_auto_in_a_valid = auto_tl_in_a_valid;
	assign fragmenter_auto_in_a_bits_opcode = auto_tl_in_a_bits_opcode;
	assign fragmenter_auto_in_a_bits_param = auto_tl_in_a_bits_param;
	assign fragmenter_auto_in_a_bits_size = auto_tl_in_a_bits_size;
	assign fragmenter_auto_in_a_bits_source = auto_tl_in_a_bits_source;
	assign fragmenter_auto_in_a_bits_address = auto_tl_in_a_bits_address;
	assign fragmenter_auto_in_a_bits_mask = auto_tl_in_a_bits_mask;
	assign fragmenter_auto_in_a_bits_data = auto_tl_in_a_bits_data;
	assign fragmenter_auto_in_a_bits_corrupt = auto_tl_in_a_bits_corrupt;
	assign fragmenter_auto_in_d_ready = auto_tl_in_d_ready;
	assign fragmenter_auto_out_a_ready = auto_control_xing_out_a_ready;
	assign fragmenter_auto_out_d_valid = auto_control_xing_out_d_valid;
	assign fragmenter_auto_out_d_bits_opcode = auto_control_xing_out_d_bits_opcode;
	assign fragmenter_auto_out_d_bits_size = auto_control_xing_out_d_bits_size;
	assign fragmenter_auto_out_d_bits_source = auto_control_xing_out_d_bits_source;
	assign fragmenter_auto_out_d_bits_data = auto_control_xing_out_d_bits_data;
endmodule
module TLMonitor_12 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [1:0] io_in_a_bits_size;
	input [7:0] io_in_a_bits_source;
	input [14:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_size;
	input [7:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_4 = io_in_a_bits_source <= 8'h9f;
	wire [4:0] _is_aligned_mask_T_1 = 5'h03 << io_in_a_bits_size;
	wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0];
	wire [14:0] _GEN_71 = {13'd0, is_aligned_mask};
	wire [14:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 15'h0000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 2'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_10 = ~_source_ok_T_4;
	wire _T_20 = io_in_a_bits_opcode == 3'h6;
	wire [14:0] _T_33 = io_in_a_bits_address ^ 15'h4000;
	wire [15:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [15:0] _T_36 = $signed(_T_34) & -16'sh1000;
	wire _T_37 = $signed(_T_36) == 16'sh0000;
	wire _T_69 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_73 = ~io_in_a_bits_mask;
	wire _T_74 = _T_73 == 4'h0;
	wire _T_78 = ~io_in_a_bits_corrupt;
	wire _T_82 = io_in_a_bits_opcode == 3'h7;
	wire _T_135 = io_in_a_bits_param != 3'h0;
	wire _T_148 = io_in_a_bits_opcode == 3'h4;
	wire _T_164 = io_in_a_bits_size <= 2'h2;
	wire _T_172 = _T_164 & _T_37;
	wire _T_183 = io_in_a_bits_param == 3'h0;
	wire _T_187 = io_in_a_bits_mask == mask;
	wire _T_195 = io_in_a_bits_opcode == 3'h0;
	wire _T_218 = _source_ok_T_4 & _T_172;
	wire _T_236 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_273 = ~mask;
	wire [3:0] _T_274 = io_in_a_bits_mask & _T_273;
	wire _T_275 = _T_274 == 4'h0;
	wire _T_279 = io_in_a_bits_opcode == 3'h2;
	wire _T_309 = io_in_a_bits_param <= 3'h4;
	wire _T_317 = io_in_a_bits_opcode == 3'h3;
	wire _T_347 = io_in_a_bits_param <= 3'h3;
	wire _T_355 = io_in_a_bits_opcode == 3'h5;
	wire _T_385 = io_in_a_bits_param <= 3'h1;
	wire _T_397 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_10 = io_in_d_bits_source <= 8'h9f;
	wire _T_401 = io_in_d_bits_opcode == 3'h6;
	wire _T_405 = io_in_d_bits_size >= 2'h2;
	wire _T_421 = io_in_d_bits_opcode == 3'h4;
	wire _T_449 = io_in_d_bits_opcode == 3'h5;
	wire _T_478 = io_in_d_bits_opcode == 3'h0;
	wire _T_495 = io_in_d_bits_opcode == 3'h1;
	wire _T_513 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [1:0] size;
	reg [7:0] source;
	reg [14:0] address;
	wire _T_543 = io_in_a_valid & ~a_first;
	wire _T_544 = io_in_a_bits_opcode == opcode;
	wire _T_548 = io_in_a_bits_param == param;
	wire _T_552 = io_in_a_bits_size == size;
	wire _T_556 = io_in_a_bits_source == source;
	wire _T_560 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] size_1;
	reg [7:0] source_1;
	wire _T_567 = io_in_d_valid & ~d_first;
	wire _T_568 = io_in_d_bits_opcode == opcode_1;
	wire _T_576 = io_in_d_bits_size == size_1;
	wire _T_580 = io_in_d_bits_source == source_1;
	reg [159:0] inflight;
	reg [639:0] inflight_opcodes;
	reg [639:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [10:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [639:0] _GEN_73 = {624'd0, _a_opcode_lookup_T_5};
	wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [639:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[639:1]};
	wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [639:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[639:1]};
	wire _T_594 = io_in_a_valid & a_first_1;
	wire [255:0] _a_set_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_a_bits_source;
	wire _T_597 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1;
	wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [10:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [2050:0] _GEN_1 = {2047'd0, a_opcodes_set_interm};
	wire [2050:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? _a_sizes_set_interm_T_1 : 3'h0);
	wire [2049:0] _GEN_2 = {2047'd0, a_sizes_set_interm};
	wire [2049:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [159:0] _T_599 = inflight >> io_in_a_bits_source;
	wire _T_601 = ~_T_599[0];
	wire [255:0] _GEN_16 = (a_first_done & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2050:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 2051'h0);
	wire [2049:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 2050'h0);
	wire _T_605 = io_in_d_valid & d_first_1;
	wire _T_607 = ~_T_401;
	wire _T_608 = (io_in_d_valid & d_first_1) & ~_T_401;
	wire [255:0] _d_clr_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_d_bits_source;
	wire [2062:0] _GEN_3 = {2047'd0, _a_opcode_lookup_T_5};
	wire [2062:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [255:0] _GEN_22 = ((d_first_done & d_first_1) & _T_607 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_23 = ((d_first_done & d_first_1) & _T_607 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_594 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [159:0] _T_618 = inflight >> io_in_d_bits_source;
	wire _T_620 = _T_618[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_625 = io_in_d_bits_opcode == _GEN_40;
	wire _T_626 = (io_in_d_bits_opcode == _GEN_32) | _T_625;
	wire _T_630 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_637 = io_in_d_bits_opcode == _GEN_56;
	wire _T_638 = (io_in_d_bits_opcode == _GEN_48) | _T_637;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {2'd0, io_in_d_bits_size};
	wire _T_642 = _GEN_82 == a_size_lookup;
	wire _T_652 = (((_T_605 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_607;
	wire _T_654 = ~io_in_d_ready | io_in_a_ready;
	wire [159:0] a_set = _GEN_16[159:0];
	wire [159:0] _inflight_T = inflight | a_set;
	wire [159:0] d_clr = _GEN_22[159:0];
	wire [159:0] _inflight_T_1 = ~d_clr;
	wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [639:0] a_opcodes_set = _GEN_19[639:0];
	wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [639:0] d_opcodes_clr = _GEN_23[639:0];
	wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [639:0] a_sizes_set = _GEN_20[639:0];
	wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_663 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [159:0] inflight_1;
	reg [639:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [639:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[639:1]};
	wire _T_689 = (io_in_d_valid & d_first_2) & _T_401;
	wire [255:0] _GEN_67 = ((d_first_done & d_first_2) & _T_401 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_68 = ((d_first_done & d_first_2) & _T_401 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire [159:0] _T_697 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_707 = _GEN_82 == c_size_lookup;
	wire [159:0] d_clr_1 = _GEN_67[159:0];
	wire [159:0] _inflight_T_4 = ~d_clr_1;
	wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0];
	wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_727 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			param <= io_in_a_bits_param;
		if (a_first_done & a_first)
			size <= io_in_a_bits_size;
		if (a_first_done & a_first)
			source <= io_in_a_bits_source;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 160'h0000000000000000000000000000000000000000;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 640'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 640'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 160'h0000000000000000000000000000000000000000;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 640'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (d_first_done)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module PeripheryBus (
	auto_coupler_to_device_named_uart_0_control_xing_out_a_ready,
	auto_coupler_to_device_named_uart_0_control_xing_out_a_valid,
	auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode,
	auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_param,
	auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size,
	auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source,
	auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address,
	auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask,
	auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data,
	auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_corrupt,
	auto_coupler_to_device_named_uart_0_control_xing_out_d_ready,
	auto_coupler_to_device_named_uart_0_control_xing_out_d_valid,
	auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode,
	auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size,
	auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source,
	auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_ready,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_valid,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_opcode,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_param,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_size,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_source,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_address,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_mask,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_data,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_corrupt,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_ready,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_valid,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_opcode,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_param,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_size,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_source,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_sink,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_denied,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_data,
	auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_corrupt,
	auto_fixedClockNode_out_clock,
	auto_fixedClockNode_out_reset,
	auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock,
	auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset,
	auto_bus_xing_in_a_ready,
	auto_bus_xing_in_a_valid,
	auto_bus_xing_in_a_bits_opcode,
	auto_bus_xing_in_a_bits_param,
	auto_bus_xing_in_a_bits_size,
	auto_bus_xing_in_a_bits_source,
	auto_bus_xing_in_a_bits_address,
	auto_bus_xing_in_a_bits_mask,
	auto_bus_xing_in_a_bits_data,
	auto_bus_xing_in_a_bits_corrupt,
	auto_bus_xing_in_d_ready,
	auto_bus_xing_in_d_valid,
	auto_bus_xing_in_d_bits_opcode,
	auto_bus_xing_in_d_bits_param,
	auto_bus_xing_in_d_bits_size,
	auto_bus_xing_in_d_bits_source,
	auto_bus_xing_in_d_bits_sink,
	auto_bus_xing_in_d_bits_denied,
	auto_bus_xing_in_d_bits_data,
	auto_bus_xing_in_d_bits_corrupt,
	clock,
	reset
);
	input auto_coupler_to_device_named_uart_0_control_xing_out_a_ready;
	output wire auto_coupler_to_device_named_uart_0_control_xing_out_a_valid;
	output wire [2:0] auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode;
	output wire [2:0] auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_param;
	output wire [1:0] auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size;
	output wire [7:0] auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source;
	output wire [30:0] auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address;
	output wire [3:0] auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask;
	output wire [31:0] auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data;
	output wire auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_corrupt;
	output wire auto_coupler_to_device_named_uart_0_control_xing_out_d_ready;
	input auto_coupler_to_device_named_uart_0_control_xing_out_d_valid;
	input [2:0] auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode;
	input [1:0] auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size;
	input [7:0] auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source;
	input [31:0] auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data;
	input auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_ready;
	output wire auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_valid;
	output wire [2:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_opcode;
	output wire [2:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_param;
	output wire [2:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_size;
	output wire [2:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_source;
	output wire [28:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_address;
	output wire [7:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_mask;
	output wire [63:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_data;
	output wire auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_corrupt;
	output wire auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_ready;
	input auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_valid;
	input [2:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_opcode;
	input [1:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_param;
	input [2:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_size;
	input [2:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_source;
	input auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_sink;
	input auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_denied;
	input [63:0] auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_data;
	input auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_corrupt;
	output wire auto_fixedClockNode_out_clock;
	output wire auto_fixedClockNode_out_reset;
	input auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock;
	input auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset;
	output wire auto_bus_xing_in_a_ready;
	input auto_bus_xing_in_a_valid;
	input [2:0] auto_bus_xing_in_a_bits_opcode;
	input [2:0] auto_bus_xing_in_a_bits_param;
	input [2:0] auto_bus_xing_in_a_bits_size;
	input [2:0] auto_bus_xing_in_a_bits_source;
	input [30:0] auto_bus_xing_in_a_bits_address;
	input [3:0] auto_bus_xing_in_a_bits_mask;
	input [31:0] auto_bus_xing_in_a_bits_data;
	input auto_bus_xing_in_a_bits_corrupt;
	input auto_bus_xing_in_d_ready;
	output wire auto_bus_xing_in_d_valid;
	output wire [2:0] auto_bus_xing_in_d_bits_opcode;
	output wire [1:0] auto_bus_xing_in_d_bits_param;
	output wire [2:0] auto_bus_xing_in_d_bits_size;
	output wire [2:0] auto_bus_xing_in_d_bits_source;
	output wire auto_bus_xing_in_d_bits_sink;
	output wire auto_bus_xing_in_d_bits_denied;
	output wire [31:0] auto_bus_xing_in_d_bits_data;
	output wire auto_bus_xing_in_d_bits_corrupt;
	output wire clock;
	output wire reset;
	wire subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_clock;
	wire subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_reset;
	wire subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_clock;
	wire subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_reset;
	wire clockGroup_auto_in_member_subsystem_pbus_0_clock;
	wire clockGroup_auto_in_member_subsystem_pbus_0_reset;
	wire clockGroup_auto_out_clock;
	wire clockGroup_auto_out_reset;
	wire fixedClockNode_auto_in_clock;
	wire fixedClockNode_auto_in_reset;
	wire fixedClockNode_auto_out_1_clock;
	wire fixedClockNode_auto_out_1_reset;
	wire fixedClockNode_auto_out_0_clock;
	wire fixedClockNode_auto_out_0_reset;
	wire fixer_clock;
	wire fixer_reset;
	wire fixer_auto_in_a_ready;
	wire fixer_auto_in_a_valid;
	wire [2:0] fixer_auto_in_a_bits_opcode;
	wire [2:0] fixer_auto_in_a_bits_param;
	wire [2:0] fixer_auto_in_a_bits_size;
	wire [2:0] fixer_auto_in_a_bits_source;
	wire [30:0] fixer_auto_in_a_bits_address;
	wire [3:0] fixer_auto_in_a_bits_mask;
	wire [31:0] fixer_auto_in_a_bits_data;
	wire fixer_auto_in_a_bits_corrupt;
	wire fixer_auto_in_d_ready;
	wire fixer_auto_in_d_valid;
	wire [2:0] fixer_auto_in_d_bits_opcode;
	wire [1:0] fixer_auto_in_d_bits_param;
	wire [2:0] fixer_auto_in_d_bits_size;
	wire [2:0] fixer_auto_in_d_bits_source;
	wire fixer_auto_in_d_bits_sink;
	wire fixer_auto_in_d_bits_denied;
	wire [31:0] fixer_auto_in_d_bits_data;
	wire fixer_auto_in_d_bits_corrupt;
	wire fixer_auto_out_a_ready;
	wire fixer_auto_out_a_valid;
	wire [2:0] fixer_auto_out_a_bits_opcode;
	wire [2:0] fixer_auto_out_a_bits_param;
	wire [2:0] fixer_auto_out_a_bits_size;
	wire [2:0] fixer_auto_out_a_bits_source;
	wire [30:0] fixer_auto_out_a_bits_address;
	wire [3:0] fixer_auto_out_a_bits_mask;
	wire [31:0] fixer_auto_out_a_bits_data;
	wire fixer_auto_out_a_bits_corrupt;
	wire fixer_auto_out_d_ready;
	wire fixer_auto_out_d_valid;
	wire [2:0] fixer_auto_out_d_bits_opcode;
	wire [1:0] fixer_auto_out_d_bits_param;
	wire [2:0] fixer_auto_out_d_bits_size;
	wire [2:0] fixer_auto_out_d_bits_source;
	wire fixer_auto_out_d_bits_sink;
	wire fixer_auto_out_d_bits_denied;
	wire [31:0] fixer_auto_out_d_bits_data;
	wire fixer_auto_out_d_bits_corrupt;
	wire in_xbar_auto_in_a_ready;
	wire in_xbar_auto_in_a_valid;
	wire [2:0] in_xbar_auto_in_a_bits_opcode;
	wire [2:0] in_xbar_auto_in_a_bits_param;
	wire [2:0] in_xbar_auto_in_a_bits_size;
	wire [2:0] in_xbar_auto_in_a_bits_source;
	wire [30:0] in_xbar_auto_in_a_bits_address;
	wire [3:0] in_xbar_auto_in_a_bits_mask;
	wire [31:0] in_xbar_auto_in_a_bits_data;
	wire in_xbar_auto_in_a_bits_corrupt;
	wire in_xbar_auto_in_d_ready;
	wire in_xbar_auto_in_d_valid;
	wire [2:0] in_xbar_auto_in_d_bits_opcode;
	wire [1:0] in_xbar_auto_in_d_bits_param;
	wire [2:0] in_xbar_auto_in_d_bits_size;
	wire [2:0] in_xbar_auto_in_d_bits_source;
	wire in_xbar_auto_in_d_bits_sink;
	wire in_xbar_auto_in_d_bits_denied;
	wire [31:0] in_xbar_auto_in_d_bits_data;
	wire in_xbar_auto_in_d_bits_corrupt;
	wire in_xbar_auto_out_a_ready;
	wire in_xbar_auto_out_a_valid;
	wire [2:0] in_xbar_auto_out_a_bits_opcode;
	wire [2:0] in_xbar_auto_out_a_bits_param;
	wire [2:0] in_xbar_auto_out_a_bits_size;
	wire [2:0] in_xbar_auto_out_a_bits_source;
	wire [30:0] in_xbar_auto_out_a_bits_address;
	wire [3:0] in_xbar_auto_out_a_bits_mask;
	wire [31:0] in_xbar_auto_out_a_bits_data;
	wire in_xbar_auto_out_a_bits_corrupt;
	wire in_xbar_auto_out_d_ready;
	wire in_xbar_auto_out_d_valid;
	wire [2:0] in_xbar_auto_out_d_bits_opcode;
	wire [1:0] in_xbar_auto_out_d_bits_param;
	wire [2:0] in_xbar_auto_out_d_bits_size;
	wire [2:0] in_xbar_auto_out_d_bits_source;
	wire in_xbar_auto_out_d_bits_sink;
	wire in_xbar_auto_out_d_bits_denied;
	wire [31:0] in_xbar_auto_out_d_bits_data;
	wire in_xbar_auto_out_d_bits_corrupt;
	wire out_xbar_clock;
	wire out_xbar_reset;
	wire out_xbar_auto_in_a_ready;
	wire out_xbar_auto_in_a_valid;
	wire [2:0] out_xbar_auto_in_a_bits_opcode;
	wire [2:0] out_xbar_auto_in_a_bits_param;
	wire [2:0] out_xbar_auto_in_a_bits_size;
	wire [2:0] out_xbar_auto_in_a_bits_source;
	wire [30:0] out_xbar_auto_in_a_bits_address;
	wire [3:0] out_xbar_auto_in_a_bits_mask;
	wire [31:0] out_xbar_auto_in_a_bits_data;
	wire out_xbar_auto_in_a_bits_corrupt;
	wire out_xbar_auto_in_d_ready;
	wire out_xbar_auto_in_d_valid;
	wire [2:0] out_xbar_auto_in_d_bits_opcode;
	wire [1:0] out_xbar_auto_in_d_bits_param;
	wire [2:0] out_xbar_auto_in_d_bits_size;
	wire [2:0] out_xbar_auto_in_d_bits_source;
	wire out_xbar_auto_in_d_bits_sink;
	wire out_xbar_auto_in_d_bits_denied;
	wire [31:0] out_xbar_auto_in_d_bits_data;
	wire out_xbar_auto_in_d_bits_corrupt;
	wire out_xbar_auto_out_2_a_ready;
	wire out_xbar_auto_out_2_a_valid;
	wire [2:0] out_xbar_auto_out_2_a_bits_opcode;
	wire [2:0] out_xbar_auto_out_2_a_bits_param;
	wire [2:0] out_xbar_auto_out_2_a_bits_size;
	wire [2:0] out_xbar_auto_out_2_a_bits_source;
	wire [30:0] out_xbar_auto_out_2_a_bits_address;
	wire [3:0] out_xbar_auto_out_2_a_bits_mask;
	wire [31:0] out_xbar_auto_out_2_a_bits_data;
	wire out_xbar_auto_out_2_a_bits_corrupt;
	wire out_xbar_auto_out_2_d_ready;
	wire out_xbar_auto_out_2_d_valid;
	wire [2:0] out_xbar_auto_out_2_d_bits_opcode;
	wire [2:0] out_xbar_auto_out_2_d_bits_size;
	wire [2:0] out_xbar_auto_out_2_d_bits_source;
	wire [31:0] out_xbar_auto_out_2_d_bits_data;
	wire out_xbar_auto_out_1_a_ready;
	wire out_xbar_auto_out_1_a_valid;
	wire [2:0] out_xbar_auto_out_1_a_bits_opcode;
	wire [2:0] out_xbar_auto_out_1_a_bits_param;
	wire [2:0] out_xbar_auto_out_1_a_bits_size;
	wire [2:0] out_xbar_auto_out_1_a_bits_source;
	wire [28:0] out_xbar_auto_out_1_a_bits_address;
	wire [3:0] out_xbar_auto_out_1_a_bits_mask;
	wire [31:0] out_xbar_auto_out_1_a_bits_data;
	wire out_xbar_auto_out_1_a_bits_corrupt;
	wire out_xbar_auto_out_1_d_ready;
	wire out_xbar_auto_out_1_d_valid;
	wire [2:0] out_xbar_auto_out_1_d_bits_opcode;
	wire [1:0] out_xbar_auto_out_1_d_bits_param;
	wire [2:0] out_xbar_auto_out_1_d_bits_size;
	wire [2:0] out_xbar_auto_out_1_d_bits_source;
	wire out_xbar_auto_out_1_d_bits_sink;
	wire out_xbar_auto_out_1_d_bits_denied;
	wire [31:0] out_xbar_auto_out_1_d_bits_data;
	wire out_xbar_auto_out_1_d_bits_corrupt;
	wire out_xbar_auto_out_0_a_ready;
	wire out_xbar_auto_out_0_a_valid;
	wire [2:0] out_xbar_auto_out_0_a_bits_opcode;
	wire [2:0] out_xbar_auto_out_0_a_bits_param;
	wire [2:0] out_xbar_auto_out_0_a_bits_size;
	wire [2:0] out_xbar_auto_out_0_a_bits_source;
	wire [14:0] out_xbar_auto_out_0_a_bits_address;
	wire [3:0] out_xbar_auto_out_0_a_bits_mask;
	wire [31:0] out_xbar_auto_out_0_a_bits_data;
	wire out_xbar_auto_out_0_a_bits_corrupt;
	wire out_xbar_auto_out_0_d_ready;
	wire out_xbar_auto_out_0_d_valid;
	wire [2:0] out_xbar_auto_out_0_d_bits_opcode;
	wire [2:0] out_xbar_auto_out_0_d_bits_size;
	wire [2:0] out_xbar_auto_out_0_d_bits_source;
	wire [31:0] out_xbar_auto_out_0_d_bits_data;
	wire buffer_clock;
	wire buffer_reset;
	wire buffer_auto_in_a_ready;
	wire buffer_auto_in_a_valid;
	wire [2:0] buffer_auto_in_a_bits_opcode;
	wire [2:0] buffer_auto_in_a_bits_param;
	wire [2:0] buffer_auto_in_a_bits_size;
	wire [2:0] buffer_auto_in_a_bits_source;
	wire [30:0] buffer_auto_in_a_bits_address;
	wire [3:0] buffer_auto_in_a_bits_mask;
	wire [31:0] buffer_auto_in_a_bits_data;
	wire buffer_auto_in_a_bits_corrupt;
	wire buffer_auto_in_d_ready;
	wire buffer_auto_in_d_valid;
	wire [2:0] buffer_auto_in_d_bits_opcode;
	wire [1:0] buffer_auto_in_d_bits_param;
	wire [2:0] buffer_auto_in_d_bits_size;
	wire [2:0] buffer_auto_in_d_bits_source;
	wire buffer_auto_in_d_bits_sink;
	wire buffer_auto_in_d_bits_denied;
	wire [31:0] buffer_auto_in_d_bits_data;
	wire buffer_auto_in_d_bits_corrupt;
	wire buffer_auto_out_a_ready;
	wire buffer_auto_out_a_valid;
	wire [2:0] buffer_auto_out_a_bits_opcode;
	wire [2:0] buffer_auto_out_a_bits_param;
	wire [2:0] buffer_auto_out_a_bits_size;
	wire [2:0] buffer_auto_out_a_bits_source;
	wire [30:0] buffer_auto_out_a_bits_address;
	wire [3:0] buffer_auto_out_a_bits_mask;
	wire [31:0] buffer_auto_out_a_bits_data;
	wire buffer_auto_out_a_bits_corrupt;
	wire buffer_auto_out_d_ready;
	wire buffer_auto_out_d_valid;
	wire [2:0] buffer_auto_out_d_bits_opcode;
	wire [1:0] buffer_auto_out_d_bits_param;
	wire [2:0] buffer_auto_out_d_bits_size;
	wire [2:0] buffer_auto_out_d_bits_source;
	wire buffer_auto_out_d_bits_sink;
	wire buffer_auto_out_d_bits_denied;
	wire [31:0] buffer_auto_out_d_bits_data;
	wire buffer_auto_out_d_bits_corrupt;
	wire atomics_clock;
	wire atomics_reset;
	wire atomics_auto_in_a_ready;
	wire atomics_auto_in_a_valid;
	wire [2:0] atomics_auto_in_a_bits_opcode;
	wire [2:0] atomics_auto_in_a_bits_param;
	wire [2:0] atomics_auto_in_a_bits_size;
	wire [2:0] atomics_auto_in_a_bits_source;
	wire [30:0] atomics_auto_in_a_bits_address;
	wire [3:0] atomics_auto_in_a_bits_mask;
	wire [31:0] atomics_auto_in_a_bits_data;
	wire atomics_auto_in_a_bits_corrupt;
	wire atomics_auto_in_d_ready;
	wire atomics_auto_in_d_valid;
	wire [2:0] atomics_auto_in_d_bits_opcode;
	wire [1:0] atomics_auto_in_d_bits_param;
	wire [2:0] atomics_auto_in_d_bits_size;
	wire [2:0] atomics_auto_in_d_bits_source;
	wire atomics_auto_in_d_bits_sink;
	wire atomics_auto_in_d_bits_denied;
	wire [31:0] atomics_auto_in_d_bits_data;
	wire atomics_auto_in_d_bits_corrupt;
	wire atomics_auto_out_a_ready;
	wire atomics_auto_out_a_valid;
	wire [2:0] atomics_auto_out_a_bits_opcode;
	wire [2:0] atomics_auto_out_a_bits_param;
	wire [2:0] atomics_auto_out_a_bits_size;
	wire [2:0] atomics_auto_out_a_bits_source;
	wire [30:0] atomics_auto_out_a_bits_address;
	wire [3:0] atomics_auto_out_a_bits_mask;
	wire [31:0] atomics_auto_out_a_bits_data;
	wire atomics_auto_out_a_bits_corrupt;
	wire atomics_auto_out_d_ready;
	wire atomics_auto_out_d_valid;
	wire [2:0] atomics_auto_out_d_bits_opcode;
	wire [1:0] atomics_auto_out_d_bits_param;
	wire [2:0] atomics_auto_out_d_bits_size;
	wire [2:0] atomics_auto_out_d_bits_source;
	wire atomics_auto_out_d_bits_sink;
	wire atomics_auto_out_d_bits_denied;
	wire [31:0] atomics_auto_out_d_bits_data;
	wire atomics_auto_out_d_bits_corrupt;
	wire buffer_1_clock;
	wire buffer_1_reset;
	wire buffer_1_auto_in_a_ready;
	wire buffer_1_auto_in_a_valid;
	wire [2:0] buffer_1_auto_in_a_bits_opcode;
	wire [2:0] buffer_1_auto_in_a_bits_param;
	wire [2:0] buffer_1_auto_in_a_bits_size;
	wire [2:0] buffer_1_auto_in_a_bits_source;
	wire [30:0] buffer_1_auto_in_a_bits_address;
	wire [3:0] buffer_1_auto_in_a_bits_mask;
	wire [31:0] buffer_1_auto_in_a_bits_data;
	wire buffer_1_auto_in_a_bits_corrupt;
	wire buffer_1_auto_in_d_ready;
	wire buffer_1_auto_in_d_valid;
	wire [2:0] buffer_1_auto_in_d_bits_opcode;
	wire [1:0] buffer_1_auto_in_d_bits_param;
	wire [2:0] buffer_1_auto_in_d_bits_size;
	wire [2:0] buffer_1_auto_in_d_bits_source;
	wire buffer_1_auto_in_d_bits_sink;
	wire buffer_1_auto_in_d_bits_denied;
	wire [31:0] buffer_1_auto_in_d_bits_data;
	wire buffer_1_auto_in_d_bits_corrupt;
	wire buffer_1_auto_out_a_ready;
	wire buffer_1_auto_out_a_valid;
	wire [2:0] buffer_1_auto_out_a_bits_opcode;
	wire [2:0] buffer_1_auto_out_a_bits_param;
	wire [2:0] buffer_1_auto_out_a_bits_size;
	wire [2:0] buffer_1_auto_out_a_bits_source;
	wire [30:0] buffer_1_auto_out_a_bits_address;
	wire [3:0] buffer_1_auto_out_a_bits_mask;
	wire [31:0] buffer_1_auto_out_a_bits_data;
	wire buffer_1_auto_out_a_bits_corrupt;
	wire buffer_1_auto_out_d_ready;
	wire buffer_1_auto_out_d_valid;
	wire [2:0] buffer_1_auto_out_d_bits_opcode;
	wire [1:0] buffer_1_auto_out_d_bits_param;
	wire [2:0] buffer_1_auto_out_d_bits_size;
	wire [2:0] buffer_1_auto_out_d_bits_source;
	wire buffer_1_auto_out_d_bits_sink;
	wire buffer_1_auto_out_d_bits_denied;
	wire [31:0] buffer_1_auto_out_d_bits_data;
	wire buffer_1_auto_out_d_bits_corrupt;
	wire coupler_to_slave_named_bootaddressreg_clock;
	wire coupler_to_slave_named_bootaddressreg_reset;
	wire coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_ready;
	wire coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_valid;
	wire [2:0] coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_opcode;
	wire [2:0] coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_param;
	wire [2:0] coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_size;
	wire [2:0] coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_source;
	wire [14:0] coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_address;
	wire [3:0] coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_mask;
	wire [31:0] coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_data;
	wire coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_corrupt;
	wire coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_ready;
	wire coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_valid;
	wire [2:0] coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_bits_opcode;
	wire [2:0] coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_bits_size;
	wire [2:0] coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_bits_source;
	wire [31:0] coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_bits_data;
	wire coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_ready;
	wire coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_valid;
	wire [2:0] coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_opcode;
	wire [2:0] coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_param;
	wire [1:0] coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_size;
	wire [7:0] coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_source;
	wire [14:0] coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_address;
	wire [3:0] coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_mask;
	wire [31:0] coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_data;
	wire coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_corrupt;
	wire coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_ready;
	wire coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_valid;
	wire [2:0] coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_bits_opcode;
	wire [1:0] coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_bits_size;
	wire [7:0] coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_bits_source;
	wire [31:0] coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_bits_data;
	wire coupler_to_port_named_serial_tl_mem_clock;
	wire coupler_to_port_named_serial_tl_mem_reset;
	wire coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_ready;
	wire coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_valid;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_opcode;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_param;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_size;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_source;
	wire [28:0] coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_address;
	wire [7:0] coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_mask;
	wire [63:0] coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_data;
	wire coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_corrupt;
	wire coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_ready;
	wire coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_valid;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_opcode;
	wire [1:0] coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_param;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_size;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_source;
	wire coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_sink;
	wire coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_denied;
	wire [63:0] coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_data;
	wire coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_corrupt;
	wire coupler_to_port_named_serial_tl_mem_auto_tl_in_a_ready;
	wire coupler_to_port_named_serial_tl_mem_auto_tl_in_a_valid;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_opcode;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_param;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_size;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_source;
	wire [28:0] coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_address;
	wire [3:0] coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_mask;
	wire [31:0] coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_data;
	wire coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_corrupt;
	wire coupler_to_port_named_serial_tl_mem_auto_tl_in_d_ready;
	wire coupler_to_port_named_serial_tl_mem_auto_tl_in_d_valid;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_opcode;
	wire [1:0] coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_param;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_size;
	wire [2:0] coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_source;
	wire coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_sink;
	wire coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_denied;
	wire [31:0] coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_data;
	wire coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_corrupt;
	wire coupler_to_device_named_uart_0_clock;
	wire coupler_to_device_named_uart_0_reset;
	wire coupler_to_device_named_uart_0_auto_control_xing_out_a_ready;
	wire coupler_to_device_named_uart_0_auto_control_xing_out_a_valid;
	wire [2:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_opcode;
	wire [2:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_param;
	wire [1:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_size;
	wire [7:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_source;
	wire [30:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_address;
	wire [3:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_mask;
	wire [31:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_data;
	wire coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_corrupt;
	wire coupler_to_device_named_uart_0_auto_control_xing_out_d_ready;
	wire coupler_to_device_named_uart_0_auto_control_xing_out_d_valid;
	wire [2:0] coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_opcode;
	wire [1:0] coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_size;
	wire [7:0] coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_source;
	wire [31:0] coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_data;
	wire coupler_to_device_named_uart_0_auto_tl_in_a_ready;
	wire coupler_to_device_named_uart_0_auto_tl_in_a_valid;
	wire [2:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_opcode;
	wire [2:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_param;
	wire [2:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_size;
	wire [2:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_source;
	wire [30:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_address;
	wire [3:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_mask;
	wire [31:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_data;
	wire coupler_to_device_named_uart_0_auto_tl_in_a_bits_corrupt;
	wire coupler_to_device_named_uart_0_auto_tl_in_d_ready;
	wire coupler_to_device_named_uart_0_auto_tl_in_d_valid;
	wire [2:0] coupler_to_device_named_uart_0_auto_tl_in_d_bits_opcode;
	wire [2:0] coupler_to_device_named_uart_0_auto_tl_in_d_bits_size;
	wire [2:0] coupler_to_device_named_uart_0_auto_tl_in_d_bits_source;
	wire [31:0] coupler_to_device_named_uart_0_auto_tl_in_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [1:0] monitor_io_in_a_bits_size;
	wire [7:0] monitor_io_in_a_bits_source;
	wire [14:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_size;
	wire [7:0] monitor_io_in_d_bits_source;
	wire bundleIn_0_clock = fixedClockNode_auto_out_0_clock;
	reg [31:0] bootAddrReg;
	wire [7:0] oldBytes_0 = bootAddrReg[7:0];
	wire [7:0] oldBytes_1 = bootAddrReg[15:8];
	wire [7:0] oldBytes_2 = bootAddrReg[23:16];
	wire [7:0] oldBytes_3 = bootAddrReg[31:24];
	wire bundleIn_0_2_a_valid = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_valid;
	wire [2:0] bundleIn_0_2_a_bits_opcode = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_opcode;
	wire in_bits_read = bundleIn_0_2_a_bits_opcode == 3'h4;
	wire [14:0] bundleIn_0_2_a_bits_address = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_address;
	wire [9:0] in_bits_index = bundleIn_0_2_a_bits_address[11:2];
	wire bundleIn_0_2_d_ready = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_ready;
	wire out_woready_0 = ((bundleIn_0_2_a_valid & bundleIn_0_2_d_ready) & ~in_bits_read) & (in_bits_index == 10'h000);
	wire [3:0] bundleIn_0_2_a_bits_mask = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_mask;
	wire [7:0] _out_backMask_T_11 = (bundleIn_0_2_a_bits_mask[3] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_9 = (bundleIn_0_2_a_bits_mask[2] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_7 = (bundleIn_0_2_a_bits_mask[1] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_5 = (bundleIn_0_2_a_bits_mask[0] ? 8'hff : 8'h00);
	wire [31:0] out_backMask = {_out_backMask_T_11, _out_backMask_T_9, _out_backMask_T_7, _out_backMask_T_5};
	wire out_womask = &out_backMask[7:0];
	wire out_f_woready = out_woready_0 & out_womask;
	wire out_womask_1 = &out_backMask[15:8];
	wire out_f_woready_1 = out_woready_0 & out_womask_1;
	wire out_womask_2 = &out_backMask[23:16];
	wire out_f_woready_2 = out_woready_0 & out_womask_2;
	wire out_womask_3 = &out_backMask[31:24];
	wire out_f_woready_3 = out_woready_0 & out_womask_3;
	wire [31:0] bundleIn_0_2_a_bits_data = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_data;
	wire [7:0] newBytes_1 = (out_f_woready_1 ? bundleIn_0_2_a_bits_data[15:8] : oldBytes_1);
	wire [7:0] newBytes_0 = (out_f_woready ? bundleIn_0_2_a_bits_data[7:0] : oldBytes_0);
	wire [7:0] newBytes_3 = (out_f_woready_3 ? bundleIn_0_2_a_bits_data[31:24] : oldBytes_3);
	wire [7:0] newBytes_2 = (out_f_woready_2 ? bundleIn_0_2_a_bits_data[23:16] : oldBytes_2);
	wire [31:0] _bootAddrReg_T = {newBytes_3, newBytes_2, newBytes_1, newBytes_0};
	wire [31:0] out_prepend_2 = {oldBytes_3, oldBytes_2, oldBytes_1, oldBytes_0};
	wire bundleIn_0_reset = fixedClockNode_auto_out_0_reset;
	ClockGroupAggregator_1 subsystem_pbus_clock_groups(
		.auto_in_member_subsystem_pbus_0_clock(subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_clock),
		.auto_in_member_subsystem_pbus_0_reset(subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_reset),
		.auto_out_member_subsystem_pbus_0_clock(subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_clock),
		.auto_out_member_subsystem_pbus_0_reset(subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_reset)
	);
	ClockGroup_1 clockGroup(
		.auto_in_member_subsystem_pbus_0_clock(clockGroup_auto_in_member_subsystem_pbus_0_clock),
		.auto_in_member_subsystem_pbus_0_reset(clockGroup_auto_in_member_subsystem_pbus_0_reset),
		.auto_out_clock(clockGroup_auto_out_clock),
		.auto_out_reset(clockGroup_auto_out_reset)
	);
	FixedClockBroadcast_1 fixedClockNode(
		.auto_in_clock(fixedClockNode_auto_in_clock),
		.auto_in_reset(fixedClockNode_auto_in_reset),
		.auto_out_1_clock(fixedClockNode_auto_out_1_clock),
		.auto_out_1_reset(fixedClockNode_auto_out_1_reset),
		.auto_out_0_clock(fixedClockNode_auto_out_0_clock),
		.auto_out_0_reset(fixedClockNode_auto_out_0_reset)
	);
	TLFIFOFixer_1 fixer(
		.clock(fixer_clock),
		.reset(fixer_reset),
		.auto_in_a_ready(fixer_auto_in_a_ready),
		.auto_in_a_valid(fixer_auto_in_a_valid),
		.auto_in_a_bits_opcode(fixer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(fixer_auto_in_a_bits_param),
		.auto_in_a_bits_size(fixer_auto_in_a_bits_size),
		.auto_in_a_bits_source(fixer_auto_in_a_bits_source),
		.auto_in_a_bits_address(fixer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(fixer_auto_in_a_bits_mask),
		.auto_in_a_bits_data(fixer_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(fixer_auto_in_a_bits_corrupt),
		.auto_in_d_ready(fixer_auto_in_d_ready),
		.auto_in_d_valid(fixer_auto_in_d_valid),
		.auto_in_d_bits_opcode(fixer_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(fixer_auto_in_d_bits_param),
		.auto_in_d_bits_size(fixer_auto_in_d_bits_size),
		.auto_in_d_bits_source(fixer_auto_in_d_bits_source),
		.auto_in_d_bits_sink(fixer_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(fixer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(fixer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(fixer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(fixer_auto_out_a_ready),
		.auto_out_a_valid(fixer_auto_out_a_valid),
		.auto_out_a_bits_opcode(fixer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(fixer_auto_out_a_bits_param),
		.auto_out_a_bits_size(fixer_auto_out_a_bits_size),
		.auto_out_a_bits_source(fixer_auto_out_a_bits_source),
		.auto_out_a_bits_address(fixer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(fixer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(fixer_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(fixer_auto_out_a_bits_corrupt),
		.auto_out_d_ready(fixer_auto_out_d_ready),
		.auto_out_d_valid(fixer_auto_out_d_valid),
		.auto_out_d_bits_opcode(fixer_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(fixer_auto_out_d_bits_param),
		.auto_out_d_bits_size(fixer_auto_out_d_bits_size),
		.auto_out_d_bits_source(fixer_auto_out_d_bits_source),
		.auto_out_d_bits_sink(fixer_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(fixer_auto_out_d_bits_denied),
		.auto_out_d_bits_data(fixer_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(fixer_auto_out_d_bits_corrupt)
	);
	TLXbar_1 in_xbar(
		.auto_in_a_ready(in_xbar_auto_in_a_ready),
		.auto_in_a_valid(in_xbar_auto_in_a_valid),
		.auto_in_a_bits_opcode(in_xbar_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(in_xbar_auto_in_a_bits_param),
		.auto_in_a_bits_size(in_xbar_auto_in_a_bits_size),
		.auto_in_a_bits_source(in_xbar_auto_in_a_bits_source),
		.auto_in_a_bits_address(in_xbar_auto_in_a_bits_address),
		.auto_in_a_bits_mask(in_xbar_auto_in_a_bits_mask),
		.auto_in_a_bits_data(in_xbar_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(in_xbar_auto_in_a_bits_corrupt),
		.auto_in_d_ready(in_xbar_auto_in_d_ready),
		.auto_in_d_valid(in_xbar_auto_in_d_valid),
		.auto_in_d_bits_opcode(in_xbar_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(in_xbar_auto_in_d_bits_param),
		.auto_in_d_bits_size(in_xbar_auto_in_d_bits_size),
		.auto_in_d_bits_source(in_xbar_auto_in_d_bits_source),
		.auto_in_d_bits_sink(in_xbar_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(in_xbar_auto_in_d_bits_denied),
		.auto_in_d_bits_data(in_xbar_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(in_xbar_auto_in_d_bits_corrupt),
		.auto_out_a_ready(in_xbar_auto_out_a_ready),
		.auto_out_a_valid(in_xbar_auto_out_a_valid),
		.auto_out_a_bits_opcode(in_xbar_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(in_xbar_auto_out_a_bits_param),
		.auto_out_a_bits_size(in_xbar_auto_out_a_bits_size),
		.auto_out_a_bits_source(in_xbar_auto_out_a_bits_source),
		.auto_out_a_bits_address(in_xbar_auto_out_a_bits_address),
		.auto_out_a_bits_mask(in_xbar_auto_out_a_bits_mask),
		.auto_out_a_bits_data(in_xbar_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(in_xbar_auto_out_a_bits_corrupt),
		.auto_out_d_ready(in_xbar_auto_out_d_ready),
		.auto_out_d_valid(in_xbar_auto_out_d_valid),
		.auto_out_d_bits_opcode(in_xbar_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(in_xbar_auto_out_d_bits_param),
		.auto_out_d_bits_size(in_xbar_auto_out_d_bits_size),
		.auto_out_d_bits_source(in_xbar_auto_out_d_bits_source),
		.auto_out_d_bits_sink(in_xbar_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(in_xbar_auto_out_d_bits_denied),
		.auto_out_d_bits_data(in_xbar_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(in_xbar_auto_out_d_bits_corrupt)
	);
	TLXbar_2 out_xbar(
		.clock(out_xbar_clock),
		.reset(out_xbar_reset),
		.auto_in_a_ready(out_xbar_auto_in_a_ready),
		.auto_in_a_valid(out_xbar_auto_in_a_valid),
		.auto_in_a_bits_opcode(out_xbar_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(out_xbar_auto_in_a_bits_param),
		.auto_in_a_bits_size(out_xbar_auto_in_a_bits_size),
		.auto_in_a_bits_source(out_xbar_auto_in_a_bits_source),
		.auto_in_a_bits_address(out_xbar_auto_in_a_bits_address),
		.auto_in_a_bits_mask(out_xbar_auto_in_a_bits_mask),
		.auto_in_a_bits_data(out_xbar_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(out_xbar_auto_in_a_bits_corrupt),
		.auto_in_d_ready(out_xbar_auto_in_d_ready),
		.auto_in_d_valid(out_xbar_auto_in_d_valid),
		.auto_in_d_bits_opcode(out_xbar_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(out_xbar_auto_in_d_bits_param),
		.auto_in_d_bits_size(out_xbar_auto_in_d_bits_size),
		.auto_in_d_bits_source(out_xbar_auto_in_d_bits_source),
		.auto_in_d_bits_sink(out_xbar_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(out_xbar_auto_in_d_bits_denied),
		.auto_in_d_bits_data(out_xbar_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(out_xbar_auto_in_d_bits_corrupt),
		.auto_out_2_a_ready(out_xbar_auto_out_2_a_ready),
		.auto_out_2_a_valid(out_xbar_auto_out_2_a_valid),
		.auto_out_2_a_bits_opcode(out_xbar_auto_out_2_a_bits_opcode),
		.auto_out_2_a_bits_param(out_xbar_auto_out_2_a_bits_param),
		.auto_out_2_a_bits_size(out_xbar_auto_out_2_a_bits_size),
		.auto_out_2_a_bits_source(out_xbar_auto_out_2_a_bits_source),
		.auto_out_2_a_bits_address(out_xbar_auto_out_2_a_bits_address),
		.auto_out_2_a_bits_mask(out_xbar_auto_out_2_a_bits_mask),
		.auto_out_2_a_bits_data(out_xbar_auto_out_2_a_bits_data),
		.auto_out_2_a_bits_corrupt(out_xbar_auto_out_2_a_bits_corrupt),
		.auto_out_2_d_ready(out_xbar_auto_out_2_d_ready),
		.auto_out_2_d_valid(out_xbar_auto_out_2_d_valid),
		.auto_out_2_d_bits_opcode(out_xbar_auto_out_2_d_bits_opcode),
		.auto_out_2_d_bits_size(out_xbar_auto_out_2_d_bits_size),
		.auto_out_2_d_bits_source(out_xbar_auto_out_2_d_bits_source),
		.auto_out_2_d_bits_data(out_xbar_auto_out_2_d_bits_data),
		.auto_out_1_a_ready(out_xbar_auto_out_1_a_ready),
		.auto_out_1_a_valid(out_xbar_auto_out_1_a_valid),
		.auto_out_1_a_bits_opcode(out_xbar_auto_out_1_a_bits_opcode),
		.auto_out_1_a_bits_param(out_xbar_auto_out_1_a_bits_param),
		.auto_out_1_a_bits_size(out_xbar_auto_out_1_a_bits_size),
		.auto_out_1_a_bits_source(out_xbar_auto_out_1_a_bits_source),
		.auto_out_1_a_bits_address(out_xbar_auto_out_1_a_bits_address),
		.auto_out_1_a_bits_mask(out_xbar_auto_out_1_a_bits_mask),
		.auto_out_1_a_bits_data(out_xbar_auto_out_1_a_bits_data),
		.auto_out_1_a_bits_corrupt(out_xbar_auto_out_1_a_bits_corrupt),
		.auto_out_1_d_ready(out_xbar_auto_out_1_d_ready),
		.auto_out_1_d_valid(out_xbar_auto_out_1_d_valid),
		.auto_out_1_d_bits_opcode(out_xbar_auto_out_1_d_bits_opcode),
		.auto_out_1_d_bits_param(out_xbar_auto_out_1_d_bits_param),
		.auto_out_1_d_bits_size(out_xbar_auto_out_1_d_bits_size),
		.auto_out_1_d_bits_source(out_xbar_auto_out_1_d_bits_source),
		.auto_out_1_d_bits_sink(out_xbar_auto_out_1_d_bits_sink),
		.auto_out_1_d_bits_denied(out_xbar_auto_out_1_d_bits_denied),
		.auto_out_1_d_bits_data(out_xbar_auto_out_1_d_bits_data),
		.auto_out_1_d_bits_corrupt(out_xbar_auto_out_1_d_bits_corrupt),
		.auto_out_0_a_ready(out_xbar_auto_out_0_a_ready),
		.auto_out_0_a_valid(out_xbar_auto_out_0_a_valid),
		.auto_out_0_a_bits_opcode(out_xbar_auto_out_0_a_bits_opcode),
		.auto_out_0_a_bits_param(out_xbar_auto_out_0_a_bits_param),
		.auto_out_0_a_bits_size(out_xbar_auto_out_0_a_bits_size),
		.auto_out_0_a_bits_source(out_xbar_auto_out_0_a_bits_source),
		.auto_out_0_a_bits_address(out_xbar_auto_out_0_a_bits_address),
		.auto_out_0_a_bits_mask(out_xbar_auto_out_0_a_bits_mask),
		.auto_out_0_a_bits_data(out_xbar_auto_out_0_a_bits_data),
		.auto_out_0_a_bits_corrupt(out_xbar_auto_out_0_a_bits_corrupt),
		.auto_out_0_d_ready(out_xbar_auto_out_0_d_ready),
		.auto_out_0_d_valid(out_xbar_auto_out_0_d_valid),
		.auto_out_0_d_bits_opcode(out_xbar_auto_out_0_d_bits_opcode),
		.auto_out_0_d_bits_size(out_xbar_auto_out_0_d_bits_size),
		.auto_out_0_d_bits_source(out_xbar_auto_out_0_d_bits_source),
		.auto_out_0_d_bits_data(out_xbar_auto_out_0_d_bits_data)
	);
	TLBuffer_1 buffer(
		.clock(buffer_clock),
		.reset(buffer_reset),
		.auto_in_a_ready(buffer_auto_in_a_ready),
		.auto_in_a_valid(buffer_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_auto_in_d_ready),
		.auto_in_d_valid(buffer_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_auto_out_a_ready),
		.auto_out_a_valid(buffer_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_auto_out_d_ready),
		.auto_out_d_valid(buffer_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(buffer_auto_out_d_bits_param),
		.auto_out_d_bits_size(buffer_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_auto_out_d_bits_source),
		.auto_out_d_bits_sink(buffer_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
		.auto_out_d_bits_data(buffer_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt)
	);
	TLAtomicAutomata atomics(
		.clock(atomics_clock),
		.reset(atomics_reset),
		.auto_in_a_ready(atomics_auto_in_a_ready),
		.auto_in_a_valid(atomics_auto_in_a_valid),
		.auto_in_a_bits_opcode(atomics_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(atomics_auto_in_a_bits_param),
		.auto_in_a_bits_size(atomics_auto_in_a_bits_size),
		.auto_in_a_bits_source(atomics_auto_in_a_bits_source),
		.auto_in_a_bits_address(atomics_auto_in_a_bits_address),
		.auto_in_a_bits_mask(atomics_auto_in_a_bits_mask),
		.auto_in_a_bits_data(atomics_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(atomics_auto_in_a_bits_corrupt),
		.auto_in_d_ready(atomics_auto_in_d_ready),
		.auto_in_d_valid(atomics_auto_in_d_valid),
		.auto_in_d_bits_opcode(atomics_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(atomics_auto_in_d_bits_param),
		.auto_in_d_bits_size(atomics_auto_in_d_bits_size),
		.auto_in_d_bits_source(atomics_auto_in_d_bits_source),
		.auto_in_d_bits_sink(atomics_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(atomics_auto_in_d_bits_denied),
		.auto_in_d_bits_data(atomics_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(atomics_auto_in_d_bits_corrupt),
		.auto_out_a_ready(atomics_auto_out_a_ready),
		.auto_out_a_valid(atomics_auto_out_a_valid),
		.auto_out_a_bits_opcode(atomics_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(atomics_auto_out_a_bits_param),
		.auto_out_a_bits_size(atomics_auto_out_a_bits_size),
		.auto_out_a_bits_source(atomics_auto_out_a_bits_source),
		.auto_out_a_bits_address(atomics_auto_out_a_bits_address),
		.auto_out_a_bits_mask(atomics_auto_out_a_bits_mask),
		.auto_out_a_bits_data(atomics_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(atomics_auto_out_a_bits_corrupt),
		.auto_out_d_ready(atomics_auto_out_d_ready),
		.auto_out_d_valid(atomics_auto_out_d_valid),
		.auto_out_d_bits_opcode(atomics_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(atomics_auto_out_d_bits_param),
		.auto_out_d_bits_size(atomics_auto_out_d_bits_size),
		.auto_out_d_bits_source(atomics_auto_out_d_bits_source),
		.auto_out_d_bits_sink(atomics_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(atomics_auto_out_d_bits_denied),
		.auto_out_d_bits_data(atomics_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(atomics_auto_out_d_bits_corrupt)
	);
	TLBuffer_2 buffer_1(
		.clock(buffer_1_clock),
		.reset(buffer_1_reset),
		.auto_in_a_ready(buffer_1_auto_in_a_ready),
		.auto_in_a_valid(buffer_1_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_1_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_1_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_1_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_1_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_1_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_1_auto_in_d_ready),
		.auto_in_d_valid(buffer_1_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_1_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_1_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_1_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_1_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_1_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_1_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_1_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_1_auto_out_a_ready),
		.auto_out_a_valid(buffer_1_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_1_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_1_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_1_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_1_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_1_auto_out_d_ready),
		.auto_out_d_valid(buffer_1_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(buffer_1_auto_out_d_bits_param),
		.auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
		.auto_out_d_bits_sink(buffer_1_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
		.auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt)
	);
	TLInterconnectCoupler_5 coupler_to_slave_named_bootaddressreg(
		.clock(coupler_to_slave_named_bootaddressreg_clock),
		.reset(coupler_to_slave_named_bootaddressreg_reset),
		.auto_buffer_in_a_ready(coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_ready),
		.auto_buffer_in_a_valid(coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_valid),
		.auto_buffer_in_a_bits_opcode(coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_opcode),
		.auto_buffer_in_a_bits_param(coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_param),
		.auto_buffer_in_a_bits_size(coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_size),
		.auto_buffer_in_a_bits_source(coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_source),
		.auto_buffer_in_a_bits_address(coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_address),
		.auto_buffer_in_a_bits_mask(coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_mask),
		.auto_buffer_in_a_bits_data(coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_data),
		.auto_buffer_in_a_bits_corrupt(coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_corrupt),
		.auto_buffer_in_d_ready(coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_ready),
		.auto_buffer_in_d_valid(coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_valid),
		.auto_buffer_in_d_bits_opcode(coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_bits_opcode),
		.auto_buffer_in_d_bits_size(coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_bits_size),
		.auto_buffer_in_d_bits_source(coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_bits_source),
		.auto_buffer_in_d_bits_data(coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_bits_data),
		.auto_fragmenter_out_a_ready(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_ready),
		.auto_fragmenter_out_a_valid(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_valid),
		.auto_fragmenter_out_a_bits_opcode(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_opcode),
		.auto_fragmenter_out_a_bits_param(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_param),
		.auto_fragmenter_out_a_bits_size(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_size),
		.auto_fragmenter_out_a_bits_source(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_source),
		.auto_fragmenter_out_a_bits_address(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_address),
		.auto_fragmenter_out_a_bits_mask(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_mask),
		.auto_fragmenter_out_a_bits_data(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_data),
		.auto_fragmenter_out_a_bits_corrupt(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_corrupt),
		.auto_fragmenter_out_d_ready(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_ready),
		.auto_fragmenter_out_d_valid(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_valid),
		.auto_fragmenter_out_d_bits_opcode(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_bits_opcode),
		.auto_fragmenter_out_d_bits_size(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_bits_size),
		.auto_fragmenter_out_d_bits_source(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_bits_source),
		.auto_fragmenter_out_d_bits_data(coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_bits_data)
	);
	TLInterconnectCoupler_6 coupler_to_port_named_serial_tl_mem(
		.clock(coupler_to_port_named_serial_tl_mem_clock),
		.reset(coupler_to_port_named_serial_tl_mem_reset),
		.auto_tlserial_manager_crossing_out_a_ready(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_ready),
		.auto_tlserial_manager_crossing_out_a_valid(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_valid),
		.auto_tlserial_manager_crossing_out_a_bits_opcode(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_opcode),
		.auto_tlserial_manager_crossing_out_a_bits_param(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_param),
		.auto_tlserial_manager_crossing_out_a_bits_size(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_size),
		.auto_tlserial_manager_crossing_out_a_bits_source(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_source),
		.auto_tlserial_manager_crossing_out_a_bits_address(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_address),
		.auto_tlserial_manager_crossing_out_a_bits_mask(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_mask),
		.auto_tlserial_manager_crossing_out_a_bits_data(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_data),
		.auto_tlserial_manager_crossing_out_a_bits_corrupt(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_corrupt),
		.auto_tlserial_manager_crossing_out_d_ready(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_ready),
		.auto_tlserial_manager_crossing_out_d_valid(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_valid),
		.auto_tlserial_manager_crossing_out_d_bits_opcode(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_opcode),
		.auto_tlserial_manager_crossing_out_d_bits_param(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_param),
		.auto_tlserial_manager_crossing_out_d_bits_size(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_size),
		.auto_tlserial_manager_crossing_out_d_bits_source(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_source),
		.auto_tlserial_manager_crossing_out_d_bits_sink(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_sink),
		.auto_tlserial_manager_crossing_out_d_bits_denied(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_denied),
		.auto_tlserial_manager_crossing_out_d_bits_data(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_data),
		.auto_tlserial_manager_crossing_out_d_bits_corrupt(coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_corrupt),
		.auto_tl_in_a_ready(coupler_to_port_named_serial_tl_mem_auto_tl_in_a_ready),
		.auto_tl_in_a_valid(coupler_to_port_named_serial_tl_mem_auto_tl_in_a_valid),
		.auto_tl_in_a_bits_opcode(coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_opcode),
		.auto_tl_in_a_bits_param(coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_param),
		.auto_tl_in_a_bits_size(coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_size),
		.auto_tl_in_a_bits_source(coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_source),
		.auto_tl_in_a_bits_address(coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_address),
		.auto_tl_in_a_bits_mask(coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_mask),
		.auto_tl_in_a_bits_data(coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_data),
		.auto_tl_in_a_bits_corrupt(coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_corrupt),
		.auto_tl_in_d_ready(coupler_to_port_named_serial_tl_mem_auto_tl_in_d_ready),
		.auto_tl_in_d_valid(coupler_to_port_named_serial_tl_mem_auto_tl_in_d_valid),
		.auto_tl_in_d_bits_opcode(coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_opcode),
		.auto_tl_in_d_bits_param(coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_param),
		.auto_tl_in_d_bits_size(coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_size),
		.auto_tl_in_d_bits_source(coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_source),
		.auto_tl_in_d_bits_sink(coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_sink),
		.auto_tl_in_d_bits_denied(coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_denied),
		.auto_tl_in_d_bits_data(coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_data),
		.auto_tl_in_d_bits_corrupt(coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_corrupt)
	);
	TLInterconnectCoupler_7 coupler_to_device_named_uart_0(
		.clock(coupler_to_device_named_uart_0_clock),
		.reset(coupler_to_device_named_uart_0_reset),
		.auto_control_xing_out_a_ready(coupler_to_device_named_uart_0_auto_control_xing_out_a_ready),
		.auto_control_xing_out_a_valid(coupler_to_device_named_uart_0_auto_control_xing_out_a_valid),
		.auto_control_xing_out_a_bits_opcode(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_opcode),
		.auto_control_xing_out_a_bits_param(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_param),
		.auto_control_xing_out_a_bits_size(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_size),
		.auto_control_xing_out_a_bits_source(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_source),
		.auto_control_xing_out_a_bits_address(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_address),
		.auto_control_xing_out_a_bits_mask(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_mask),
		.auto_control_xing_out_a_bits_data(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_data),
		.auto_control_xing_out_a_bits_corrupt(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_corrupt),
		.auto_control_xing_out_d_ready(coupler_to_device_named_uart_0_auto_control_xing_out_d_ready),
		.auto_control_xing_out_d_valid(coupler_to_device_named_uart_0_auto_control_xing_out_d_valid),
		.auto_control_xing_out_d_bits_opcode(coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_opcode),
		.auto_control_xing_out_d_bits_size(coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_size),
		.auto_control_xing_out_d_bits_source(coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_source),
		.auto_control_xing_out_d_bits_data(coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_data),
		.auto_tl_in_a_ready(coupler_to_device_named_uart_0_auto_tl_in_a_ready),
		.auto_tl_in_a_valid(coupler_to_device_named_uart_0_auto_tl_in_a_valid),
		.auto_tl_in_a_bits_opcode(coupler_to_device_named_uart_0_auto_tl_in_a_bits_opcode),
		.auto_tl_in_a_bits_param(coupler_to_device_named_uart_0_auto_tl_in_a_bits_param),
		.auto_tl_in_a_bits_size(coupler_to_device_named_uart_0_auto_tl_in_a_bits_size),
		.auto_tl_in_a_bits_source(coupler_to_device_named_uart_0_auto_tl_in_a_bits_source),
		.auto_tl_in_a_bits_address(coupler_to_device_named_uart_0_auto_tl_in_a_bits_address),
		.auto_tl_in_a_bits_mask(coupler_to_device_named_uart_0_auto_tl_in_a_bits_mask),
		.auto_tl_in_a_bits_data(coupler_to_device_named_uart_0_auto_tl_in_a_bits_data),
		.auto_tl_in_a_bits_corrupt(coupler_to_device_named_uart_0_auto_tl_in_a_bits_corrupt),
		.auto_tl_in_d_ready(coupler_to_device_named_uart_0_auto_tl_in_d_ready),
		.auto_tl_in_d_valid(coupler_to_device_named_uart_0_auto_tl_in_d_valid),
		.auto_tl_in_d_bits_opcode(coupler_to_device_named_uart_0_auto_tl_in_d_bits_opcode),
		.auto_tl_in_d_bits_size(coupler_to_device_named_uart_0_auto_tl_in_d_bits_size),
		.auto_tl_in_d_bits_source(coupler_to_device_named_uart_0_auto_tl_in_d_bits_source),
		.auto_tl_in_d_bits_data(coupler_to_device_named_uart_0_auto_tl_in_d_bits_data)
	);
	TLMonitor_12 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	assign auto_coupler_to_device_named_uart_0_control_xing_out_a_valid = coupler_to_device_named_uart_0_auto_control_xing_out_a_valid;
	assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode = coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_opcode;
	assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_param = coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_param;
	assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size = coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_size;
	assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source = coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_source;
	assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address = coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_address;
	assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask = coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_mask;
	assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data = coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_data;
	assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_corrupt = coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_corrupt;
	assign auto_coupler_to_device_named_uart_0_control_xing_out_d_ready = coupler_to_device_named_uart_0_auto_control_xing_out_d_ready;
	assign auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_valid = coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_valid;
	assign auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_opcode = coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_opcode;
	assign auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_param = coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_param;
	assign auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_size = coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_size;
	assign auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_source = coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_source;
	assign auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_address = coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_address;
	assign auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_mask = coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_mask;
	assign auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_data = coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_data;
	assign auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_corrupt = coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_bits_corrupt;
	assign auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_ready = coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_ready;
	assign auto_fixedClockNode_out_clock = fixedClockNode_auto_out_1_clock;
	assign auto_fixedClockNode_out_reset = fixedClockNode_auto_out_1_reset;
	assign auto_bus_xing_in_a_ready = buffer_1_auto_in_a_ready;
	assign auto_bus_xing_in_d_valid = buffer_1_auto_in_d_valid;
	assign auto_bus_xing_in_d_bits_opcode = buffer_1_auto_in_d_bits_opcode;
	assign auto_bus_xing_in_d_bits_param = buffer_1_auto_in_d_bits_param;
	assign auto_bus_xing_in_d_bits_size = buffer_1_auto_in_d_bits_size;
	assign auto_bus_xing_in_d_bits_source = buffer_1_auto_in_d_bits_source;
	assign auto_bus_xing_in_d_bits_sink = buffer_1_auto_in_d_bits_sink;
	assign auto_bus_xing_in_d_bits_denied = buffer_1_auto_in_d_bits_denied;
	assign auto_bus_xing_in_d_bits_data = buffer_1_auto_in_d_bits_data;
	assign auto_bus_xing_in_d_bits_corrupt = buffer_1_auto_in_d_bits_corrupt;
	assign clock = fixedClockNode_auto_out_0_clock;
	assign reset = fixedClockNode_auto_out_0_reset;
	assign subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_clock = auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock;
	assign subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_reset = auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset;
	assign clockGroup_auto_in_member_subsystem_pbus_0_clock = subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_clock;
	assign clockGroup_auto_in_member_subsystem_pbus_0_reset = subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_reset;
	assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock;
	assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset;
	assign fixer_clock = fixedClockNode_auto_out_0_clock;
	assign fixer_reset = fixedClockNode_auto_out_0_reset;
	assign fixer_auto_in_a_valid = buffer_auto_out_a_valid;
	assign fixer_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode;
	assign fixer_auto_in_a_bits_param = buffer_auto_out_a_bits_param;
	assign fixer_auto_in_a_bits_size = buffer_auto_out_a_bits_size;
	assign fixer_auto_in_a_bits_source = buffer_auto_out_a_bits_source;
	assign fixer_auto_in_a_bits_address = buffer_auto_out_a_bits_address;
	assign fixer_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask;
	assign fixer_auto_in_a_bits_data = buffer_auto_out_a_bits_data;
	assign fixer_auto_in_a_bits_corrupt = buffer_auto_out_a_bits_corrupt;
	assign fixer_auto_in_d_ready = buffer_auto_out_d_ready;
	assign fixer_auto_out_a_ready = out_xbar_auto_in_a_ready;
	assign fixer_auto_out_d_valid = out_xbar_auto_in_d_valid;
	assign fixer_auto_out_d_bits_opcode = out_xbar_auto_in_d_bits_opcode;
	assign fixer_auto_out_d_bits_param = out_xbar_auto_in_d_bits_param;
	assign fixer_auto_out_d_bits_size = out_xbar_auto_in_d_bits_size;
	assign fixer_auto_out_d_bits_source = out_xbar_auto_in_d_bits_source;
	assign fixer_auto_out_d_bits_sink = out_xbar_auto_in_d_bits_sink;
	assign fixer_auto_out_d_bits_denied = out_xbar_auto_in_d_bits_denied;
	assign fixer_auto_out_d_bits_data = out_xbar_auto_in_d_bits_data;
	assign fixer_auto_out_d_bits_corrupt = out_xbar_auto_in_d_bits_corrupt;
	assign in_xbar_auto_in_a_valid = buffer_1_auto_out_a_valid;
	assign in_xbar_auto_in_a_bits_opcode = buffer_1_auto_out_a_bits_opcode;
	assign in_xbar_auto_in_a_bits_param = buffer_1_auto_out_a_bits_param;
	assign in_xbar_auto_in_a_bits_size = buffer_1_auto_out_a_bits_size;
	assign in_xbar_auto_in_a_bits_source = buffer_1_auto_out_a_bits_source;
	assign in_xbar_auto_in_a_bits_address = buffer_1_auto_out_a_bits_address;
	assign in_xbar_auto_in_a_bits_mask = buffer_1_auto_out_a_bits_mask;
	assign in_xbar_auto_in_a_bits_data = buffer_1_auto_out_a_bits_data;
	assign in_xbar_auto_in_a_bits_corrupt = buffer_1_auto_out_a_bits_corrupt;
	assign in_xbar_auto_in_d_ready = buffer_1_auto_out_d_ready;
	assign in_xbar_auto_out_a_ready = atomics_auto_in_a_ready;
	assign in_xbar_auto_out_d_valid = atomics_auto_in_d_valid;
	assign in_xbar_auto_out_d_bits_opcode = atomics_auto_in_d_bits_opcode;
	assign in_xbar_auto_out_d_bits_param = atomics_auto_in_d_bits_param;
	assign in_xbar_auto_out_d_bits_size = atomics_auto_in_d_bits_size;
	assign in_xbar_auto_out_d_bits_source = atomics_auto_in_d_bits_source;
	assign in_xbar_auto_out_d_bits_sink = atomics_auto_in_d_bits_sink;
	assign in_xbar_auto_out_d_bits_denied = atomics_auto_in_d_bits_denied;
	assign in_xbar_auto_out_d_bits_data = atomics_auto_in_d_bits_data;
	assign in_xbar_auto_out_d_bits_corrupt = atomics_auto_in_d_bits_corrupt;
	assign out_xbar_clock = fixedClockNode_auto_out_0_clock;
	assign out_xbar_reset = fixedClockNode_auto_out_0_reset;
	assign out_xbar_auto_in_a_valid = fixer_auto_out_a_valid;
	assign out_xbar_auto_in_a_bits_opcode = fixer_auto_out_a_bits_opcode;
	assign out_xbar_auto_in_a_bits_param = fixer_auto_out_a_bits_param;
	assign out_xbar_auto_in_a_bits_size = fixer_auto_out_a_bits_size;
	assign out_xbar_auto_in_a_bits_source = fixer_auto_out_a_bits_source;
	assign out_xbar_auto_in_a_bits_address = fixer_auto_out_a_bits_address;
	assign out_xbar_auto_in_a_bits_mask = fixer_auto_out_a_bits_mask;
	assign out_xbar_auto_in_a_bits_data = fixer_auto_out_a_bits_data;
	assign out_xbar_auto_in_a_bits_corrupt = fixer_auto_out_a_bits_corrupt;
	assign out_xbar_auto_in_d_ready = fixer_auto_out_d_ready;
	assign out_xbar_auto_out_2_a_ready = coupler_to_device_named_uart_0_auto_tl_in_a_ready;
	assign out_xbar_auto_out_2_d_valid = coupler_to_device_named_uart_0_auto_tl_in_d_valid;
	assign out_xbar_auto_out_2_d_bits_opcode = coupler_to_device_named_uart_0_auto_tl_in_d_bits_opcode;
	assign out_xbar_auto_out_2_d_bits_size = coupler_to_device_named_uart_0_auto_tl_in_d_bits_size;
	assign out_xbar_auto_out_2_d_bits_source = coupler_to_device_named_uart_0_auto_tl_in_d_bits_source;
	assign out_xbar_auto_out_2_d_bits_data = coupler_to_device_named_uart_0_auto_tl_in_d_bits_data;
	assign out_xbar_auto_out_1_a_ready = coupler_to_port_named_serial_tl_mem_auto_tl_in_a_ready;
	assign out_xbar_auto_out_1_d_valid = coupler_to_port_named_serial_tl_mem_auto_tl_in_d_valid;
	assign out_xbar_auto_out_1_d_bits_opcode = coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_opcode;
	assign out_xbar_auto_out_1_d_bits_param = coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_param;
	assign out_xbar_auto_out_1_d_bits_size = coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_size;
	assign out_xbar_auto_out_1_d_bits_source = coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_source;
	assign out_xbar_auto_out_1_d_bits_sink = coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_sink;
	assign out_xbar_auto_out_1_d_bits_denied = coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_denied;
	assign out_xbar_auto_out_1_d_bits_data = coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_data;
	assign out_xbar_auto_out_1_d_bits_corrupt = coupler_to_port_named_serial_tl_mem_auto_tl_in_d_bits_corrupt;
	assign out_xbar_auto_out_0_a_ready = coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_ready;
	assign out_xbar_auto_out_0_d_valid = coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_valid;
	assign out_xbar_auto_out_0_d_bits_opcode = coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_bits_opcode;
	assign out_xbar_auto_out_0_d_bits_size = coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_bits_size;
	assign out_xbar_auto_out_0_d_bits_source = coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_bits_source;
	assign out_xbar_auto_out_0_d_bits_data = coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_bits_data;
	assign buffer_clock = fixedClockNode_auto_out_0_clock;
	assign buffer_reset = fixedClockNode_auto_out_0_reset;
	assign buffer_auto_in_a_valid = atomics_auto_out_a_valid;
	assign buffer_auto_in_a_bits_opcode = atomics_auto_out_a_bits_opcode;
	assign buffer_auto_in_a_bits_param = atomics_auto_out_a_bits_param;
	assign buffer_auto_in_a_bits_size = atomics_auto_out_a_bits_size;
	assign buffer_auto_in_a_bits_source = atomics_auto_out_a_bits_source;
	assign buffer_auto_in_a_bits_address = atomics_auto_out_a_bits_address;
	assign buffer_auto_in_a_bits_mask = atomics_auto_out_a_bits_mask;
	assign buffer_auto_in_a_bits_data = atomics_auto_out_a_bits_data;
	assign buffer_auto_in_a_bits_corrupt = atomics_auto_out_a_bits_corrupt;
	assign buffer_auto_in_d_ready = atomics_auto_out_d_ready;
	assign buffer_auto_out_a_ready = fixer_auto_in_a_ready;
	assign buffer_auto_out_d_valid = fixer_auto_in_d_valid;
	assign buffer_auto_out_d_bits_opcode = fixer_auto_in_d_bits_opcode;
	assign buffer_auto_out_d_bits_param = fixer_auto_in_d_bits_param;
	assign buffer_auto_out_d_bits_size = fixer_auto_in_d_bits_size;
	assign buffer_auto_out_d_bits_source = fixer_auto_in_d_bits_source;
	assign buffer_auto_out_d_bits_sink = fixer_auto_in_d_bits_sink;
	assign buffer_auto_out_d_bits_denied = fixer_auto_in_d_bits_denied;
	assign buffer_auto_out_d_bits_data = fixer_auto_in_d_bits_data;
	assign buffer_auto_out_d_bits_corrupt = fixer_auto_in_d_bits_corrupt;
	assign atomics_clock = fixedClockNode_auto_out_0_clock;
	assign atomics_reset = fixedClockNode_auto_out_0_reset;
	assign atomics_auto_in_a_valid = in_xbar_auto_out_a_valid;
	assign atomics_auto_in_a_bits_opcode = in_xbar_auto_out_a_bits_opcode;
	assign atomics_auto_in_a_bits_param = in_xbar_auto_out_a_bits_param;
	assign atomics_auto_in_a_bits_size = in_xbar_auto_out_a_bits_size;
	assign atomics_auto_in_a_bits_source = in_xbar_auto_out_a_bits_source;
	assign atomics_auto_in_a_bits_address = in_xbar_auto_out_a_bits_address;
	assign atomics_auto_in_a_bits_mask = in_xbar_auto_out_a_bits_mask;
	assign atomics_auto_in_a_bits_data = in_xbar_auto_out_a_bits_data;
	assign atomics_auto_in_a_bits_corrupt = in_xbar_auto_out_a_bits_corrupt;
	assign atomics_auto_in_d_ready = in_xbar_auto_out_d_ready;
	assign atomics_auto_out_a_ready = buffer_auto_in_a_ready;
	assign atomics_auto_out_d_valid = buffer_auto_in_d_valid;
	assign atomics_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode;
	assign atomics_auto_out_d_bits_param = buffer_auto_in_d_bits_param;
	assign atomics_auto_out_d_bits_size = buffer_auto_in_d_bits_size;
	assign atomics_auto_out_d_bits_source = buffer_auto_in_d_bits_source;
	assign atomics_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink;
	assign atomics_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied;
	assign atomics_auto_out_d_bits_data = buffer_auto_in_d_bits_data;
	assign atomics_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt;
	assign buffer_1_clock = fixedClockNode_auto_out_0_clock;
	assign buffer_1_reset = fixedClockNode_auto_out_0_reset;
	assign buffer_1_auto_in_a_valid = auto_bus_xing_in_a_valid;
	assign buffer_1_auto_in_a_bits_opcode = auto_bus_xing_in_a_bits_opcode;
	assign buffer_1_auto_in_a_bits_param = auto_bus_xing_in_a_bits_param;
	assign buffer_1_auto_in_a_bits_size = auto_bus_xing_in_a_bits_size;
	assign buffer_1_auto_in_a_bits_source = auto_bus_xing_in_a_bits_source;
	assign buffer_1_auto_in_a_bits_address = auto_bus_xing_in_a_bits_address;
	assign buffer_1_auto_in_a_bits_mask = auto_bus_xing_in_a_bits_mask;
	assign buffer_1_auto_in_a_bits_data = auto_bus_xing_in_a_bits_data;
	assign buffer_1_auto_in_a_bits_corrupt = auto_bus_xing_in_a_bits_corrupt;
	assign buffer_1_auto_in_d_ready = auto_bus_xing_in_d_ready;
	assign buffer_1_auto_out_a_ready = in_xbar_auto_in_a_ready;
	assign buffer_1_auto_out_d_valid = in_xbar_auto_in_d_valid;
	assign buffer_1_auto_out_d_bits_opcode = in_xbar_auto_in_d_bits_opcode;
	assign buffer_1_auto_out_d_bits_param = in_xbar_auto_in_d_bits_param;
	assign buffer_1_auto_out_d_bits_size = in_xbar_auto_in_d_bits_size;
	assign buffer_1_auto_out_d_bits_source = in_xbar_auto_in_d_bits_source;
	assign buffer_1_auto_out_d_bits_sink = in_xbar_auto_in_d_bits_sink;
	assign buffer_1_auto_out_d_bits_denied = in_xbar_auto_in_d_bits_denied;
	assign buffer_1_auto_out_d_bits_data = in_xbar_auto_in_d_bits_data;
	assign buffer_1_auto_out_d_bits_corrupt = in_xbar_auto_in_d_bits_corrupt;
	assign coupler_to_slave_named_bootaddressreg_clock = fixedClockNode_auto_out_0_clock;
	assign coupler_to_slave_named_bootaddressreg_reset = fixedClockNode_auto_out_0_reset;
	assign coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_valid = out_xbar_auto_out_0_a_valid;
	assign coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_opcode = out_xbar_auto_out_0_a_bits_opcode;
	assign coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_param = out_xbar_auto_out_0_a_bits_param;
	assign coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_size = out_xbar_auto_out_0_a_bits_size;
	assign coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_source = out_xbar_auto_out_0_a_bits_source;
	assign coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_address = out_xbar_auto_out_0_a_bits_address;
	assign coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_mask = out_xbar_auto_out_0_a_bits_mask;
	assign coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_data = out_xbar_auto_out_0_a_bits_data;
	assign coupler_to_slave_named_bootaddressreg_auto_buffer_in_a_bits_corrupt = out_xbar_auto_out_0_a_bits_corrupt;
	assign coupler_to_slave_named_bootaddressreg_auto_buffer_in_d_ready = out_xbar_auto_out_0_d_ready;
	assign coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_ready = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_ready;
	assign coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_valid = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_valid;
	assign coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_bits_opcode = {2'd0, in_bits_read};
	assign coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_bits_size = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_size;
	assign coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_bits_source = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_source;
	assign coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_bits_data = (in_bits_index == 10'h000 ? out_prepend_2 : 32'h00000000);
	assign coupler_to_port_named_serial_tl_mem_clock = fixedClockNode_auto_out_0_clock;
	assign coupler_to_port_named_serial_tl_mem_reset = fixedClockNode_auto_out_0_reset;
	assign coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_a_ready = auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_ready;
	assign coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_valid = auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_valid;
	assign coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_opcode = auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_opcode;
	assign coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_param = auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_param;
	assign coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_size = auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_size;
	assign coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_source = auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_source;
	assign coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_sink = auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_sink;
	assign coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_denied = auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_denied;
	assign coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_data = auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_data;
	assign coupler_to_port_named_serial_tl_mem_auto_tlserial_manager_crossing_out_d_bits_corrupt = auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_corrupt;
	assign coupler_to_port_named_serial_tl_mem_auto_tl_in_a_valid = out_xbar_auto_out_1_a_valid;
	assign coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_opcode = out_xbar_auto_out_1_a_bits_opcode;
	assign coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_param = out_xbar_auto_out_1_a_bits_param;
	assign coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_size = out_xbar_auto_out_1_a_bits_size;
	assign coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_source = out_xbar_auto_out_1_a_bits_source;
	assign coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_address = out_xbar_auto_out_1_a_bits_address;
	assign coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_mask = out_xbar_auto_out_1_a_bits_mask;
	assign coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_data = out_xbar_auto_out_1_a_bits_data;
	assign coupler_to_port_named_serial_tl_mem_auto_tl_in_a_bits_corrupt = out_xbar_auto_out_1_a_bits_corrupt;
	assign coupler_to_port_named_serial_tl_mem_auto_tl_in_d_ready = out_xbar_auto_out_1_d_ready;
	assign coupler_to_device_named_uart_0_clock = fixedClockNode_auto_out_0_clock;
	assign coupler_to_device_named_uart_0_reset = fixedClockNode_auto_out_0_reset;
	assign coupler_to_device_named_uart_0_auto_control_xing_out_a_ready = auto_coupler_to_device_named_uart_0_control_xing_out_a_ready;
	assign coupler_to_device_named_uart_0_auto_control_xing_out_d_valid = auto_coupler_to_device_named_uart_0_control_xing_out_d_valid;
	assign coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_opcode = auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode;
	assign coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_size = auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size;
	assign coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_source = auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source;
	assign coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_data = auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data;
	assign coupler_to_device_named_uart_0_auto_tl_in_a_valid = out_xbar_auto_out_2_a_valid;
	assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_opcode = out_xbar_auto_out_2_a_bits_opcode;
	assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_param = out_xbar_auto_out_2_a_bits_param;
	assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_size = out_xbar_auto_out_2_a_bits_size;
	assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_source = out_xbar_auto_out_2_a_bits_source;
	assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_address = out_xbar_auto_out_2_a_bits_address;
	assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_mask = out_xbar_auto_out_2_a_bits_mask;
	assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_data = out_xbar_auto_out_2_a_bits_data;
	assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_corrupt = out_xbar_auto_out_2_a_bits_corrupt;
	assign coupler_to_device_named_uart_0_auto_tl_in_d_ready = out_xbar_auto_out_2_d_ready;
	assign monitor_clock = fixedClockNode_auto_out_0_clock;
	assign monitor_reset = fixedClockNode_auto_out_0_reset;
	assign monitor_io_in_a_ready = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_ready;
	assign monitor_io_in_a_valid = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_valid;
	assign monitor_io_in_a_bits_opcode = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_opcode;
	assign monitor_io_in_a_bits_param = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_param;
	assign monitor_io_in_a_bits_size = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_size;
	assign monitor_io_in_a_bits_source = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_source;
	assign monitor_io_in_a_bits_address = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_address;
	assign monitor_io_in_a_bits_mask = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_corrupt;
	assign monitor_io_in_d_ready = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_d_ready;
	assign monitor_io_in_d_valid = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_valid;
	assign monitor_io_in_d_bits_opcode = {2'd0, in_bits_read};
	assign monitor_io_in_d_bits_size = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_size;
	assign monitor_io_in_d_bits_source = coupler_to_slave_named_bootaddressreg_auto_fragmenter_out_a_bits_source;
	always @(posedge bundleIn_0_clock)
		if (bundleIn_0_reset)
			bootAddrReg <= 32'h80000000;
		else if (((out_f_woready | out_f_woready_1) | out_f_woready_2) | out_f_woready_3)
			bootAddrReg <= _bootAddrReg_T;
endmodule
module ClockGroupAggregator_2 (
	auto_in_member_subsystem_fbus_0_clock,
	auto_in_member_subsystem_fbus_0_reset,
	auto_out_member_subsystem_fbus_0_clock,
	auto_out_member_subsystem_fbus_0_reset
);
	input auto_in_member_subsystem_fbus_0_clock;
	input auto_in_member_subsystem_fbus_0_reset;
	output wire auto_out_member_subsystem_fbus_0_clock;
	output wire auto_out_member_subsystem_fbus_0_reset;
	assign auto_out_member_subsystem_fbus_0_clock = auto_in_member_subsystem_fbus_0_clock;
	assign auto_out_member_subsystem_fbus_0_reset = auto_in_member_subsystem_fbus_0_reset;
endmodule
module ClockGroup_2 (
	auto_in_member_subsystem_fbus_0_clock,
	auto_in_member_subsystem_fbus_0_reset,
	auto_out_clock,
	auto_out_reset
);
	input auto_in_member_subsystem_fbus_0_clock;
	input auto_in_member_subsystem_fbus_0_reset;
	output wire auto_out_clock;
	output wire auto_out_reset;
	assign auto_out_clock = auto_in_member_subsystem_fbus_0_clock;
	assign auto_out_reset = auto_in_member_subsystem_fbus_0_reset;
endmodule
module TLXbar_3 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module TLMonitor_13 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = ~io_in_a_bits_source;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_5 = ~_source_ok_T;
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_15 = io_in_a_bits_opcode == 3'h6;
	wire _T_17 = io_in_a_bits_size <= 4'hc;
	wire _T_20 = _T_17 & _source_ok_T;
	wire [32:0] _T_26 = $signed(_T_7) & -33'sh000005000;
	wire _T_27 = $signed(_T_26) == 33'sh000000000;
	wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_29 = {1'b0, $signed(_T_28)};
	wire [32:0] _T_31 = $signed(_T_29) & -33'sh000001000;
	wire _T_32 = $signed(_T_31) == 33'sh000000000;
	wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [32:0] _T_36 = $signed(_T_34) & -33'sh000010000;
	wire _T_37 = $signed(_T_36) == 33'sh000000000;
	wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_39 = {1'b0, $signed(_T_38)};
	wire [32:0] _T_41 = $signed(_T_39) & -33'sh000010000;
	wire _T_42 = $signed(_T_41) == 33'sh000000000;
	wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_44 = {1'b0, $signed(_T_43)};
	wire [32:0] _T_46 = $signed(_T_44) & -33'sh000011000;
	wire _T_47 = $signed(_T_46) == 33'sh000000000;
	wire [31:0] _T_48 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_49 = {1'b0, $signed(_T_48)};
	wire [32:0] _T_51 = $signed(_T_49) & -33'sh000010000;
	wire _T_52 = $signed(_T_51) == 33'sh000000000;
	wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_54 = {1'b0, $signed(_T_53)};
	wire [32:0] _T_56 = $signed(_T_54) & -33'sh004000000;
	wire _T_57 = $signed(_T_56) == 33'sh000000000;
	wire [31:0] _T_58 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_59 = {1'b0, $signed(_T_58)};
	wire [32:0] _T_61 = $signed(_T_59) & -33'sh000001000;
	wire _T_62 = $signed(_T_61) == 33'sh000000000;
	wire [31:0] _T_63 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_64 = {1'b0, $signed(_T_63)};
	wire [32:0] _T_66 = $signed(_T_64) & -33'sh000001000;
	wire _T_67 = $signed(_T_66) == 33'sh000000000;
	wire [31:0] _T_68 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_69 = {1'b0, $signed(_T_68)};
	wire [32:0] _T_71 = $signed(_T_69) & -33'sh000004000;
	wire _T_72 = $signed(_T_71) == 33'sh000000000;
	wire _T_167 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_171 = ~io_in_a_bits_mask;
	wire _T_172 = _T_171 == 4'h0;
	wire _T_176 = ~io_in_a_bits_corrupt;
	wire _T_180 = io_in_a_bits_opcode == 3'h7;
	wire _T_336 = io_in_a_bits_param != 3'h0;
	wire _T_349 = io_in_a_bits_opcode == 3'h4;
	wire _T_368 = _T_17 & _T_32;
	wire _T_370 = io_in_a_bits_size <= 4'h6;
	wire _T_425 = (((((((_T_27 | _T_37) | _T_42) | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_426 = _T_370 & _T_425;
	wire _T_428 = _T_368 | _T_426;
	wire _T_438 = io_in_a_bits_param == 3'h0;
	wire _T_442 = io_in_a_bits_mask == mask;
	wire _T_450 = io_in_a_bits_opcode == 3'h0;
	wire _T_511 = (((((_T_27 | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_512 = _T_370 & _T_511;
	wire _T_527 = _T_368 | _T_512;
	wire _T_529 = _T_20 & _T_527;
	wire _T_547 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_640 = ~mask;
	wire [3:0] _T_641 = io_in_a_bits_mask & _T_640;
	wire _T_642 = _T_641 == 4'h0;
	wire _T_646 = io_in_a_bits_opcode == 3'h2;
	wire _T_654 = io_in_a_bits_size <= 4'h2;
	wire _T_703 = ((((((_T_27 | _T_32) | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_704 = _T_654 & _T_703;
	wire _T_720 = _T_20 & _T_704;
	wire _T_730 = io_in_a_bits_param <= 3'h4;
	wire _T_738 = io_in_a_bits_opcode == 3'h3;
	wire _T_822 = io_in_a_bits_param <= 3'h3;
	wire _T_830 = io_in_a_bits_opcode == 3'h5;
	wire _T_904 = _T_20 & _T_368;
	wire _T_914 = io_in_a_bits_param <= 3'h1;
	wire _T_926 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_1 = ~io_in_d_bits_source;
	wire _T_930 = io_in_d_bits_opcode == 3'h6;
	wire _T_934 = io_in_d_bits_size >= 4'h2;
	wire _T_938 = io_in_d_bits_param == 2'h0;
	wire _T_942 = ~io_in_d_bits_corrupt;
	wire _T_946 = ~io_in_d_bits_denied;
	wire _T_950 = io_in_d_bits_opcode == 3'h4;
	wire _T_961 = io_in_d_bits_param <= 2'h2;
	wire _T_965 = io_in_d_bits_param != 2'h2;
	wire _T_978 = io_in_d_bits_opcode == 3'h5;
	wire _T_998 = _T_946 | io_in_d_bits_corrupt;
	wire _T_1007 = io_in_d_bits_opcode == 3'h0;
	wire _T_1024 = io_in_d_bits_opcode == 3'h1;
	wire _T_1042 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg source;
	reg [31:0] address;
	wire _T_1072 = io_in_a_valid & ~a_first;
	wire _T_1073 = io_in_a_bits_opcode == opcode;
	wire _T_1077 = io_in_a_bits_param == param;
	wire _T_1081 = io_in_a_bits_size == size;
	wire _T_1085 = io_in_a_bits_source == source;
	wire _T_1089 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg source_1;
	reg sink;
	reg denied;
	wire _T_1096 = io_in_d_valid & ~d_first;
	wire _T_1097 = io_in_d_bits_opcode == opcode_1;
	wire _T_1101 = io_in_d_bits_param == param_1;
	wire _T_1105 = io_in_d_bits_size == size_1;
	wire _T_1109 = io_in_d_bits_source == source_1;
	wire _T_1113 = io_in_d_bits_sink == sink;
	wire _T_1117 = io_in_d_bits_denied == denied;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [7:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [3:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_73 = {12'd0, _a_opcode_lookup_T_1};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0};
	wire [7:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T;
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [15:0] _GEN_75 = {8'd0, _a_size_lookup_T_1};
	wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_size_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_1123 = io_in_a_valid & a_first_1;
	wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source;
	wire [1:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire _T_1126 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [2:0] _GEN_77 = {io_in_a_bits_source, 2'h0};
	wire [3:0] _a_opcodes_set_T = {1'd0, _GEN_77};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _GEN_1 = {15'd0, a_opcodes_set_interm};
	wire [18:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [19:0] _GEN_2 = {15'd0, a_sizes_set_interm};
	wire [19:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire _T_1130 = ~(inflight >> io_in_a_bits_source);
	wire [1:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire [18:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [19:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 20'h00000);
	wire _T_1134 = io_in_d_valid & d_first_1;
	wire _T_1136 = ~_T_930;
	wire _T_1137 = (io_in_d_valid & d_first_1) & ~_T_930;
	wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source;
	wire [1:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_930 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_3 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [30:0] _GEN_4 = {15'd0, _a_size_lookup_T_5};
	wire [30:0] _d_sizes_clr_T_5 = _GEN_4 << _a_size_lookup_T;
	wire [1:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_1136 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1136 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [30:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1136 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_1123 & (io_in_a_bits_source == io_in_d_bits_source);
	wire _T_1149 = (inflight >> io_in_d_bits_source) | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1154 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1155 = (io_in_d_bits_opcode == _GEN_32) | _T_1154;
	wire _T_1159 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1166 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1167 = (io_in_d_bits_opcode == _GEN_48) | _T_1166;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_79 = {4'd0, io_in_d_bits_size};
	wire _T_1171 = _GEN_79 == a_size_lookup;
	wire _T_1181 = (((_T_1134 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_1136;
	wire _T_1183 = ~io_in_d_ready | io_in_a_ready;
	wire a_set_wo_ready = _GEN_15[0];
	wire d_clr_wo_ready = _GEN_21[0];
	wire _T_1190 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire a_set = _GEN_16[0];
	wire d_clr = _GEN_22[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [7:0] a_sizes_set = _GEN_20[7:0];
	wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [7:0] d_sizes_clr = _GEN_24[7:0];
	wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1199 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [7:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [7:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T;
	wire [15:0] _GEN_83 = {8'd0, _c_size_lookup_T_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_83 & _a_size_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_1225 = (io_in_d_valid & d_first_2) & _T_930;
	wire [30:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_930 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire _T_1233 = 1'h0 >> io_in_d_bits_source;
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1243 = _GEN_79 == c_size_lookup;
	wire [7:0] d_sizes_clr_1 = _GEN_69[7:0];
	wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 8'h00;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 8'h00;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module Queue_4 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_data,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [3:0] io_enq_bits_size;
	input io_enq_bits_source;
	input [31:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input [31:0] io_enq_bits_data;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [3:0] io_deq_bits_size;
	output wire io_deq_bits_source;
	output wire [31:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire [31:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg [2:0] ram_opcode [0:1];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [2:0] ram_param [0:1];
	wire ram_param_io_deq_bits_MPORT_en;
	wire ram_param_io_deq_bits_MPORT_addr;
	wire [2:0] ram_param_io_deq_bits_MPORT_data;
	wire [2:0] ram_param_MPORT_data;
	wire ram_param_MPORT_addr;
	wire ram_param_MPORT_mask;
	wire ram_param_MPORT_en;
	reg [3:0] ram_size [0:1];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [3:0] ram_size_io_deq_bits_MPORT_data;
	wire [3:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg ram_source [0:1];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire ram_source_io_deq_bits_MPORT_data;
	wire ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg [31:0] ram_address [0:1];
	wire ram_address_io_deq_bits_MPORT_en;
	wire ram_address_io_deq_bits_MPORT_addr;
	wire [31:0] ram_address_io_deq_bits_MPORT_data;
	wire [31:0] ram_address_MPORT_data;
	wire ram_address_MPORT_addr;
	wire ram_address_MPORT_mask;
	wire ram_address_MPORT_en;
	reg [3:0] ram_mask [0:1];
	wire ram_mask_io_deq_bits_MPORT_en;
	wire ram_mask_io_deq_bits_MPORT_addr;
	wire [3:0] ram_mask_io_deq_bits_MPORT_data;
	wire [3:0] ram_mask_MPORT_data;
	wire ram_mask_MPORT_addr;
	wire ram_mask_MPORT_mask;
	wire ram_mask_MPORT_en;
	reg [31:0] ram_data [0:1];
	wire ram_data_io_deq_bits_MPORT_en;
	wire ram_data_io_deq_bits_MPORT_addr;
	wire [31:0] ram_data_io_deq_bits_MPORT_data;
	wire [31:0] ram_data_MPORT_data;
	wire ram_data_MPORT_addr;
	wire ram_data_MPORT_mask;
	wire ram_data_MPORT_en;
	reg ram_corrupt [0:1];
	wire ram_corrupt_io_deq_bits_MPORT_en;
	wire ram_corrupt_io_deq_bits_MPORT_addr;
	wire ram_corrupt_io_deq_bits_MPORT_data;
	wire ram_corrupt_MPORT_data;
	wire ram_corrupt_MPORT_addr;
	wire ram_corrupt_MPORT_mask;
	wire ram_corrupt_MPORT_en;
	reg value;
	reg value_1;
	reg maybe_full;
	wire ptr_match = value == value_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = value;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_param_io_deq_bits_MPORT_en = 1'h1;
	assign ram_param_io_deq_bits_MPORT_addr = value_1;
	assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr];
	assign ram_param_MPORT_data = io_enq_bits_param;
	assign ram_param_MPORT_addr = value;
	assign ram_param_MPORT_mask = 1'h1;
	assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = value_1;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = value;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = value_1;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = value;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_address_io_deq_bits_MPORT_en = 1'h1;
	assign ram_address_io_deq_bits_MPORT_addr = value_1;
	assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr];
	assign ram_address_MPORT_data = io_enq_bits_address;
	assign ram_address_MPORT_addr = value;
	assign ram_address_MPORT_mask = 1'h1;
	assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
	assign ram_mask_io_deq_bits_MPORT_addr = value_1;
	assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr];
	assign ram_mask_MPORT_data = io_enq_bits_mask;
	assign ram_mask_MPORT_addr = value;
	assign ram_mask_MPORT_mask = 1'h1;
	assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_data_io_deq_bits_MPORT_en = 1'h1;
	assign ram_data_io_deq_bits_MPORT_addr = value_1;
	assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr];
	assign ram_data_MPORT_data = io_enq_bits_data;
	assign ram_data_MPORT_addr = value;
	assign ram_data_MPORT_mask = 1'h1;
	assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
	assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
	assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr];
	assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
	assign ram_corrupt_MPORT_addr = value;
	assign ram_corrupt_MPORT_mask = 1'h1;
	assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data;
	assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data;
	assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data;
	assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_param_MPORT_en & ram_param_MPORT_mask)
			ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (ram_address_MPORT_en & ram_address_MPORT_mask)
			ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data;
		if (ram_mask_MPORT_en & ram_mask_MPORT_mask)
			ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data;
		if (ram_data_MPORT_en & ram_data_MPORT_mask)
			ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data;
		if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask)
			ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data;
		if (reset)
			value <= 1'h0;
		else if (do_enq)
			value <= value + 1'h1;
		if (reset)
			value_1 <= 1'h0;
		else if (do_deq)
			value_1 <= value_1 + 1'h1;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module Queue_5 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_sink,
	io_enq_bits_denied,
	io_enq_bits_data,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_sink,
	io_deq_bits_denied,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [1:0] io_enq_bits_param;
	input [3:0] io_enq_bits_size;
	input io_enq_bits_source;
	input io_enq_bits_sink;
	input io_enq_bits_denied;
	input [31:0] io_enq_bits_data;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [1:0] io_deq_bits_param;
	output wire [3:0] io_deq_bits_size;
	output wire io_deq_bits_source;
	output wire io_deq_bits_sink;
	output wire io_deq_bits_denied;
	output wire [31:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg [2:0] ram_opcode [0:1];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [1:0] ram_param [0:1];
	wire ram_param_io_deq_bits_MPORT_en;
	wire ram_param_io_deq_bits_MPORT_addr;
	wire [1:0] ram_param_io_deq_bits_MPORT_data;
	wire [1:0] ram_param_MPORT_data;
	wire ram_param_MPORT_addr;
	wire ram_param_MPORT_mask;
	wire ram_param_MPORT_en;
	reg [3:0] ram_size [0:1];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [3:0] ram_size_io_deq_bits_MPORT_data;
	wire [3:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg ram_source [0:1];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire ram_source_io_deq_bits_MPORT_data;
	wire ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg ram_sink [0:1];
	wire ram_sink_io_deq_bits_MPORT_en;
	wire ram_sink_io_deq_bits_MPORT_addr;
	wire ram_sink_io_deq_bits_MPORT_data;
	wire ram_sink_MPORT_data;
	wire ram_sink_MPORT_addr;
	wire ram_sink_MPORT_mask;
	wire ram_sink_MPORT_en;
	reg ram_denied [0:1];
	wire ram_denied_io_deq_bits_MPORT_en;
	wire ram_denied_io_deq_bits_MPORT_addr;
	wire ram_denied_io_deq_bits_MPORT_data;
	wire ram_denied_MPORT_data;
	wire ram_denied_MPORT_addr;
	wire ram_denied_MPORT_mask;
	wire ram_denied_MPORT_en;
	reg [31:0] ram_data [0:1];
	wire ram_data_io_deq_bits_MPORT_en;
	wire ram_data_io_deq_bits_MPORT_addr;
	wire [31:0] ram_data_io_deq_bits_MPORT_data;
	wire [31:0] ram_data_MPORT_data;
	wire ram_data_MPORT_addr;
	wire ram_data_MPORT_mask;
	wire ram_data_MPORT_en;
	reg ram_corrupt [0:1];
	wire ram_corrupt_io_deq_bits_MPORT_en;
	wire ram_corrupt_io_deq_bits_MPORT_addr;
	wire ram_corrupt_io_deq_bits_MPORT_data;
	wire ram_corrupt_MPORT_data;
	wire ram_corrupt_MPORT_addr;
	wire ram_corrupt_MPORT_mask;
	wire ram_corrupt_MPORT_en;
	reg value;
	reg value_1;
	reg maybe_full;
	wire ptr_match = value == value_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = value;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_param_io_deq_bits_MPORT_en = 1'h1;
	assign ram_param_io_deq_bits_MPORT_addr = value_1;
	assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr];
	assign ram_param_MPORT_data = io_enq_bits_param;
	assign ram_param_MPORT_addr = value;
	assign ram_param_MPORT_mask = 1'h1;
	assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = value_1;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = value;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = value_1;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = value;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_sink_io_deq_bits_MPORT_en = 1'h1;
	assign ram_sink_io_deq_bits_MPORT_addr = value_1;
	assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr];
	assign ram_sink_MPORT_data = io_enq_bits_sink;
	assign ram_sink_MPORT_addr = value;
	assign ram_sink_MPORT_mask = 1'h1;
	assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_denied_io_deq_bits_MPORT_en = 1'h1;
	assign ram_denied_io_deq_bits_MPORT_addr = value_1;
	assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr];
	assign ram_denied_MPORT_data = io_enq_bits_denied;
	assign ram_denied_MPORT_addr = value;
	assign ram_denied_MPORT_mask = 1'h1;
	assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_data_io_deq_bits_MPORT_en = 1'h1;
	assign ram_data_io_deq_bits_MPORT_addr = value_1;
	assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr];
	assign ram_data_MPORT_data = io_enq_bits_data;
	assign ram_data_MPORT_addr = value;
	assign ram_data_MPORT_mask = 1'h1;
	assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
	assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
	assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr];
	assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
	assign ram_corrupt_MPORT_addr = value;
	assign ram_corrupt_MPORT_mask = 1'h1;
	assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data;
	assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data;
	assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data;
	assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_param_MPORT_en & ram_param_MPORT_mask)
			ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (ram_sink_MPORT_en & ram_sink_MPORT_mask)
			ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data;
		if (ram_denied_MPORT_en & ram_denied_MPORT_mask)
			ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data;
		if (ram_data_MPORT_en & ram_data_MPORT_mask)
			ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data;
		if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask)
			ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data;
		if (reset)
			value <= 1'h0;
		else if (do_enq)
			value <= value + 1'h1;
		if (reset)
			value_1 <= 1'h0;
		else if (do_deq)
			value_1 <= value_1 + 1'h1;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module TLBuffer_4 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire monitor_io_in_a_bits_source;
	wire [31:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [3:0] monitor_io_in_d_bits_size;
	wire monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire bundleOut_0_a_q_clock;
	wire bundleOut_0_a_q_reset;
	wire bundleOut_0_a_q_io_enq_ready;
	wire bundleOut_0_a_q_io_enq_valid;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_param;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_size;
	wire bundleOut_0_a_q_io_enq_bits_source;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_data;
	wire bundleOut_0_a_q_io_enq_bits_corrupt;
	wire bundleOut_0_a_q_io_deq_ready;
	wire bundleOut_0_a_q_io_deq_valid;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_param;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_size;
	wire bundleOut_0_a_q_io_deq_bits_source;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_data;
	wire bundleOut_0_a_q_io_deq_bits_corrupt;
	wire bundleIn_0_d_q_clock;
	wire bundleIn_0_d_q_reset;
	wire bundleIn_0_d_q_io_enq_ready;
	wire bundleIn_0_d_q_io_enq_valid;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_enq_bits_param;
	wire [3:0] bundleIn_0_d_q_io_enq_bits_size;
	wire bundleIn_0_d_q_io_enq_bits_source;
	wire bundleIn_0_d_q_io_enq_bits_sink;
	wire bundleIn_0_d_q_io_enq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_enq_bits_data;
	wire bundleIn_0_d_q_io_enq_bits_corrupt;
	wire bundleIn_0_d_q_io_deq_ready;
	wire bundleIn_0_d_q_io_deq_valid;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_param;
	wire [3:0] bundleIn_0_d_q_io_deq_bits_size;
	wire bundleIn_0_d_q_io_deq_bits_source;
	wire bundleIn_0_d_q_io_deq_bits_sink;
	wire bundleIn_0_d_q_io_deq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_deq_bits_data;
	wire bundleIn_0_d_q_io_deq_bits_corrupt;
	TLMonitor_13 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Queue_4 bundleOut_0_a_q(
		.clock(bundleOut_0_a_q_clock),
		.reset(bundleOut_0_a_q_reset),
		.io_enq_ready(bundleOut_0_a_q_io_enq_ready),
		.io_enq_valid(bundleOut_0_a_q_io_enq_valid),
		.io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
		.io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
		.io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
		.io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
		.io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
		.io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleOut_0_a_q_io_deq_ready),
		.io_deq_valid(bundleOut_0_a_q_io_deq_valid),
		.io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
		.io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
		.io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
		.io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
		.io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
		.io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
	);
	Queue_5 bundleIn_0_d_q(
		.clock(bundleIn_0_d_q_clock),
		.reset(bundleIn_0_d_q_reset),
		.io_enq_ready(bundleIn_0_d_q_io_enq_ready),
		.io_enq_valid(bundleIn_0_d_q_io_enq_valid),
		.io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
		.io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
		.io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
		.io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
		.io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
		.io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleIn_0_d_q_io_deq_ready),
		.io_deq_valid(bundleIn_0_d_q_io_deq_valid),
		.io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
		.io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
		.io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
		.io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
		.io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
		.io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data;
	assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid;
	assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode;
	assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param;
	assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size;
	assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source;
	assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address;
	assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask;
	assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data;
	assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt;
	assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign bundleOut_0_a_q_clock = clock;
	assign bundleOut_0_a_q_reset = reset;
	assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid;
	assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param;
	assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size;
	assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source;
	assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address;
	assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask;
	assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data;
	assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready;
	assign bundleIn_0_d_q_clock = clock;
	assign bundleIn_0_d_q_reset = reset;
	assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid;
	assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign bundleIn_0_d_q_io_enq_bits_param = auto_out_d_bits_param;
	assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size;
	assign bundleIn_0_d_q_io_enq_bits_source = 1'h0;
	assign bundleIn_0_d_q_io_enq_bits_sink = auto_out_d_bits_sink;
	assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied;
	assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data;
	assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt;
	assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready;
endmodule
module TLMonitor_14 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = ~io_in_a_bits_source;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_5 = ~_source_ok_T;
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_15 = io_in_a_bits_opcode == 3'h6;
	wire _T_17 = io_in_a_bits_size <= 4'hc;
	wire _T_20 = _T_17 & _source_ok_T;
	wire [32:0] _T_26 = $signed(_T_7) & -33'sh000005000;
	wire _T_27 = $signed(_T_26) == 33'sh000000000;
	wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_29 = {1'b0, $signed(_T_28)};
	wire [32:0] _T_31 = $signed(_T_29) & -33'sh000001000;
	wire _T_32 = $signed(_T_31) == 33'sh000000000;
	wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [32:0] _T_36 = $signed(_T_34) & -33'sh000010000;
	wire _T_37 = $signed(_T_36) == 33'sh000000000;
	wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_39 = {1'b0, $signed(_T_38)};
	wire [32:0] _T_41 = $signed(_T_39) & -33'sh000010000;
	wire _T_42 = $signed(_T_41) == 33'sh000000000;
	wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_44 = {1'b0, $signed(_T_43)};
	wire [32:0] _T_46 = $signed(_T_44) & -33'sh000011000;
	wire _T_47 = $signed(_T_46) == 33'sh000000000;
	wire [31:0] _T_48 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_49 = {1'b0, $signed(_T_48)};
	wire [32:0] _T_51 = $signed(_T_49) & -33'sh000010000;
	wire _T_52 = $signed(_T_51) == 33'sh000000000;
	wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_54 = {1'b0, $signed(_T_53)};
	wire [32:0] _T_56 = $signed(_T_54) & -33'sh004000000;
	wire _T_57 = $signed(_T_56) == 33'sh000000000;
	wire [31:0] _T_58 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_59 = {1'b0, $signed(_T_58)};
	wire [32:0] _T_61 = $signed(_T_59) & -33'sh000001000;
	wire _T_62 = $signed(_T_61) == 33'sh000000000;
	wire [31:0] _T_63 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_64 = {1'b0, $signed(_T_63)};
	wire [32:0] _T_66 = $signed(_T_64) & -33'sh000001000;
	wire _T_67 = $signed(_T_66) == 33'sh000000000;
	wire [31:0] _T_68 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_69 = {1'b0, $signed(_T_68)};
	wire [32:0] _T_71 = $signed(_T_69) & -33'sh000004000;
	wire _T_72 = $signed(_T_71) == 33'sh000000000;
	wire _T_167 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_171 = ~io_in_a_bits_mask;
	wire _T_172 = _T_171 == 4'h0;
	wire _T_176 = ~io_in_a_bits_corrupt;
	wire _T_180 = io_in_a_bits_opcode == 3'h7;
	wire _T_336 = io_in_a_bits_param != 3'h0;
	wire _T_349 = io_in_a_bits_opcode == 3'h4;
	wire _T_368 = _T_17 & _T_32;
	wire _T_370 = io_in_a_bits_size <= 4'h6;
	wire _T_425 = (((((((_T_27 | _T_37) | _T_42) | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_426 = _T_370 & _T_425;
	wire _T_428 = _T_368 | _T_426;
	wire _T_438 = io_in_a_bits_param == 3'h0;
	wire _T_442 = io_in_a_bits_mask == mask;
	wire _T_450 = io_in_a_bits_opcode == 3'h0;
	wire _T_511 = (((((_T_27 | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_512 = _T_370 & _T_511;
	wire _T_527 = _T_368 | _T_512;
	wire _T_529 = _T_20 & _T_527;
	wire _T_547 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_640 = ~mask;
	wire [3:0] _T_641 = io_in_a_bits_mask & _T_640;
	wire _T_642 = _T_641 == 4'h0;
	wire _T_646 = io_in_a_bits_opcode == 3'h2;
	wire _T_654 = io_in_a_bits_size <= 4'h2;
	wire _T_703 = ((((((_T_27 | _T_32) | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_704 = _T_654 & _T_703;
	wire _T_720 = _T_20 & _T_704;
	wire _T_730 = io_in_a_bits_param <= 3'h4;
	wire _T_738 = io_in_a_bits_opcode == 3'h3;
	wire _T_822 = io_in_a_bits_param <= 3'h3;
	wire _T_830 = io_in_a_bits_opcode == 3'h5;
	wire _T_904 = _T_20 & _T_368;
	wire _T_914 = io_in_a_bits_param <= 3'h1;
	wire _T_926 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_1 = ~io_in_d_bits_source;
	wire _T_930 = io_in_d_bits_opcode == 3'h6;
	wire _T_934 = io_in_d_bits_size >= 4'h2;
	wire _T_938 = io_in_d_bits_param == 2'h0;
	wire _T_942 = ~io_in_d_bits_corrupt;
	wire _T_946 = ~io_in_d_bits_denied;
	wire _T_950 = io_in_d_bits_opcode == 3'h4;
	wire _T_961 = io_in_d_bits_param <= 2'h2;
	wire _T_965 = io_in_d_bits_param != 2'h2;
	wire _T_978 = io_in_d_bits_opcode == 3'h5;
	wire _T_998 = _T_946 | io_in_d_bits_corrupt;
	wire _T_1007 = io_in_d_bits_opcode == 3'h0;
	wire _T_1024 = io_in_d_bits_opcode == 3'h1;
	wire _T_1042 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg source;
	reg [31:0] address;
	wire _T_1072 = io_in_a_valid & ~a_first;
	wire _T_1073 = io_in_a_bits_opcode == opcode;
	wire _T_1077 = io_in_a_bits_param == param;
	wire _T_1081 = io_in_a_bits_size == size;
	wire _T_1085 = io_in_a_bits_source == source;
	wire _T_1089 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg source_1;
	reg sink;
	reg denied;
	wire _T_1096 = io_in_d_valid & ~d_first;
	wire _T_1097 = io_in_d_bits_opcode == opcode_1;
	wire _T_1101 = io_in_d_bits_param == param_1;
	wire _T_1105 = io_in_d_bits_size == size_1;
	wire _T_1109 = io_in_d_bits_source == source_1;
	wire _T_1113 = io_in_d_bits_sink == sink;
	wire _T_1117 = io_in_d_bits_denied == denied;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [7:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [3:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_73 = {12'd0, _a_opcode_lookup_T_1};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0};
	wire [7:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T;
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [15:0] _GEN_75 = {8'd0, _a_size_lookup_T_1};
	wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_size_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_1123 = io_in_a_valid & a_first_1;
	wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source;
	wire [1:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire _T_1126 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [2:0] _GEN_77 = {io_in_a_bits_source, 2'h0};
	wire [3:0] _a_opcodes_set_T = {1'd0, _GEN_77};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _GEN_1 = {15'd0, a_opcodes_set_interm};
	wire [18:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [19:0] _GEN_2 = {15'd0, a_sizes_set_interm};
	wire [19:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire _T_1130 = ~(inflight >> io_in_a_bits_source);
	wire [1:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire [18:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [19:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 20'h00000);
	wire _T_1134 = io_in_d_valid & d_first_1;
	wire _T_1136 = ~_T_930;
	wire _T_1137 = (io_in_d_valid & d_first_1) & ~_T_930;
	wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source;
	wire [1:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_930 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_3 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [30:0] _GEN_4 = {15'd0, _a_size_lookup_T_5};
	wire [30:0] _d_sizes_clr_T_5 = _GEN_4 << _a_size_lookup_T;
	wire [1:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_1136 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1136 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [30:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1136 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_1123 & (io_in_a_bits_source == io_in_d_bits_source);
	wire _T_1149 = (inflight >> io_in_d_bits_source) | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1154 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1155 = (io_in_d_bits_opcode == _GEN_32) | _T_1154;
	wire _T_1159 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1166 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1167 = (io_in_d_bits_opcode == _GEN_48) | _T_1166;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_79 = {4'd0, io_in_d_bits_size};
	wire _T_1171 = _GEN_79 == a_size_lookup;
	wire _T_1181 = (((_T_1134 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_1136;
	wire _T_1183 = ~io_in_d_ready | io_in_a_ready;
	wire a_set_wo_ready = _GEN_15[0];
	wire d_clr_wo_ready = _GEN_21[0];
	wire _T_1190 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire a_set = _GEN_16[0];
	wire d_clr = _GEN_22[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [7:0] a_sizes_set = _GEN_20[7:0];
	wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [7:0] d_sizes_clr = _GEN_24[7:0];
	wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1199 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [7:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [7:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T;
	wire [15:0] _GEN_83 = {8'd0, _c_size_lookup_T_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_83 & _a_size_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_1225 = (io_in_d_valid & d_first_2) & _T_930;
	wire [30:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_930 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire _T_1233 = 1'h0 >> io_in_d_bits_source;
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1243 = _GEN_79 == c_size_lookup;
	wire [7:0] d_sizes_clr_1 = _GEN_69[7:0];
	wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 8'h00;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 8'h00;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module TLBuffer_5 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire monitor_io_in_a_bits_source;
	wire [31:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [3:0] monitor_io_in_d_bits_size;
	wire monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire bundleOut_0_a_q_clock;
	wire bundleOut_0_a_q_reset;
	wire bundleOut_0_a_q_io_enq_ready;
	wire bundleOut_0_a_q_io_enq_valid;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_param;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_size;
	wire bundleOut_0_a_q_io_enq_bits_source;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_data;
	wire bundleOut_0_a_q_io_enq_bits_corrupt;
	wire bundleOut_0_a_q_io_deq_ready;
	wire bundleOut_0_a_q_io_deq_valid;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_param;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_size;
	wire bundleOut_0_a_q_io_deq_bits_source;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_data;
	wire bundleOut_0_a_q_io_deq_bits_corrupt;
	wire bundleIn_0_d_q_clock;
	wire bundleIn_0_d_q_reset;
	wire bundleIn_0_d_q_io_enq_ready;
	wire bundleIn_0_d_q_io_enq_valid;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_enq_bits_param;
	wire [3:0] bundleIn_0_d_q_io_enq_bits_size;
	wire bundleIn_0_d_q_io_enq_bits_source;
	wire bundleIn_0_d_q_io_enq_bits_sink;
	wire bundleIn_0_d_q_io_enq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_enq_bits_data;
	wire bundleIn_0_d_q_io_enq_bits_corrupt;
	wire bundleIn_0_d_q_io_deq_ready;
	wire bundleIn_0_d_q_io_deq_valid;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_param;
	wire [3:0] bundleIn_0_d_q_io_deq_bits_size;
	wire bundleIn_0_d_q_io_deq_bits_source;
	wire bundleIn_0_d_q_io_deq_bits_sink;
	wire bundleIn_0_d_q_io_deq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_deq_bits_data;
	wire bundleIn_0_d_q_io_deq_bits_corrupt;
	TLMonitor_14 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Queue_4 bundleOut_0_a_q(
		.clock(bundleOut_0_a_q_clock),
		.reset(bundleOut_0_a_q_reset),
		.io_enq_ready(bundleOut_0_a_q_io_enq_ready),
		.io_enq_valid(bundleOut_0_a_q_io_enq_valid),
		.io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
		.io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
		.io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
		.io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
		.io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
		.io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleOut_0_a_q_io_deq_ready),
		.io_deq_valid(bundleOut_0_a_q_io_deq_valid),
		.io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
		.io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
		.io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
		.io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
		.io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
		.io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
	);
	Queue_5 bundleIn_0_d_q(
		.clock(bundleIn_0_d_q_clock),
		.reset(bundleIn_0_d_q_reset),
		.io_enq_ready(bundleIn_0_d_q_io_enq_ready),
		.io_enq_valid(bundleIn_0_d_q_io_enq_valid),
		.io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
		.io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
		.io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
		.io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
		.io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
		.io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleIn_0_d_q_io_deq_ready),
		.io_deq_valid(bundleIn_0_d_q_io_deq_valid),
		.io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
		.io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
		.io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
		.io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
		.io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
		.io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data;
	assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid;
	assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode;
	assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param;
	assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size;
	assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source;
	assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address;
	assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask;
	assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data;
	assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt;
	assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign bundleOut_0_a_q_clock = clock;
	assign bundleOut_0_a_q_reset = reset;
	assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid;
	assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param;
	assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size;
	assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source;
	assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address;
	assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask;
	assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data;
	assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready;
	assign bundleIn_0_d_q_clock = clock;
	assign bundleIn_0_d_q_reset = reset;
	assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid;
	assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign bundleIn_0_d_q_io_enq_bits_param = auto_out_d_bits_param;
	assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size;
	assign bundleIn_0_d_q_io_enq_bits_source = 1'h0;
	assign bundleIn_0_d_q_io_enq_bits_sink = auto_out_d_bits_sink;
	assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied;
	assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data;
	assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt;
	assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready;
endmodule
module TLInterconnectCoupler_8 (
	clock,
	reset,
	auto_buffer_in_a_ready,
	auto_buffer_in_a_valid,
	auto_buffer_in_a_bits_opcode,
	auto_buffer_in_a_bits_param,
	auto_buffer_in_a_bits_size,
	auto_buffer_in_a_bits_source,
	auto_buffer_in_a_bits_address,
	auto_buffer_in_a_bits_mask,
	auto_buffer_in_a_bits_data,
	auto_buffer_in_a_bits_corrupt,
	auto_buffer_in_d_ready,
	auto_buffer_in_d_valid,
	auto_buffer_in_d_bits_opcode,
	auto_buffer_in_d_bits_param,
	auto_buffer_in_d_bits_size,
	auto_buffer_in_d_bits_source,
	auto_buffer_in_d_bits_sink,
	auto_buffer_in_d_bits_denied,
	auto_buffer_in_d_bits_data,
	auto_buffer_in_d_bits_corrupt,
	auto_tl_out_a_ready,
	auto_tl_out_a_valid,
	auto_tl_out_a_bits_opcode,
	auto_tl_out_a_bits_param,
	auto_tl_out_a_bits_size,
	auto_tl_out_a_bits_source,
	auto_tl_out_a_bits_address,
	auto_tl_out_a_bits_mask,
	auto_tl_out_a_bits_data,
	auto_tl_out_a_bits_corrupt,
	auto_tl_out_d_ready,
	auto_tl_out_d_valid,
	auto_tl_out_d_bits_opcode,
	auto_tl_out_d_bits_param,
	auto_tl_out_d_bits_size,
	auto_tl_out_d_bits_sink,
	auto_tl_out_d_bits_denied,
	auto_tl_out_d_bits_data,
	auto_tl_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_buffer_in_a_ready;
	input auto_buffer_in_a_valid;
	input [2:0] auto_buffer_in_a_bits_opcode;
	input [2:0] auto_buffer_in_a_bits_param;
	input [3:0] auto_buffer_in_a_bits_size;
	input auto_buffer_in_a_bits_source;
	input [31:0] auto_buffer_in_a_bits_address;
	input [3:0] auto_buffer_in_a_bits_mask;
	input [31:0] auto_buffer_in_a_bits_data;
	input auto_buffer_in_a_bits_corrupt;
	input auto_buffer_in_d_ready;
	output wire auto_buffer_in_d_valid;
	output wire [2:0] auto_buffer_in_d_bits_opcode;
	output wire [1:0] auto_buffer_in_d_bits_param;
	output wire [3:0] auto_buffer_in_d_bits_size;
	output wire auto_buffer_in_d_bits_source;
	output wire auto_buffer_in_d_bits_sink;
	output wire auto_buffer_in_d_bits_denied;
	output wire [31:0] auto_buffer_in_d_bits_data;
	output wire auto_buffer_in_d_bits_corrupt;
	input auto_tl_out_a_ready;
	output wire auto_tl_out_a_valid;
	output wire [2:0] auto_tl_out_a_bits_opcode;
	output wire [2:0] auto_tl_out_a_bits_param;
	output wire [3:0] auto_tl_out_a_bits_size;
	output wire auto_tl_out_a_bits_source;
	output wire [31:0] auto_tl_out_a_bits_address;
	output wire [3:0] auto_tl_out_a_bits_mask;
	output wire [31:0] auto_tl_out_a_bits_data;
	output wire auto_tl_out_a_bits_corrupt;
	output wire auto_tl_out_d_ready;
	input auto_tl_out_d_valid;
	input [2:0] auto_tl_out_d_bits_opcode;
	input [1:0] auto_tl_out_d_bits_param;
	input [3:0] auto_tl_out_d_bits_size;
	input auto_tl_out_d_bits_sink;
	input auto_tl_out_d_bits_denied;
	input [31:0] auto_tl_out_d_bits_data;
	input auto_tl_out_d_bits_corrupt;
	wire buffer_clock;
	wire buffer_reset;
	wire buffer_auto_in_a_ready;
	wire buffer_auto_in_a_valid;
	wire [2:0] buffer_auto_in_a_bits_opcode;
	wire [2:0] buffer_auto_in_a_bits_param;
	wire [3:0] buffer_auto_in_a_bits_size;
	wire buffer_auto_in_a_bits_source;
	wire [31:0] buffer_auto_in_a_bits_address;
	wire [3:0] buffer_auto_in_a_bits_mask;
	wire [31:0] buffer_auto_in_a_bits_data;
	wire buffer_auto_in_a_bits_corrupt;
	wire buffer_auto_in_d_ready;
	wire buffer_auto_in_d_valid;
	wire [2:0] buffer_auto_in_d_bits_opcode;
	wire [1:0] buffer_auto_in_d_bits_param;
	wire [3:0] buffer_auto_in_d_bits_size;
	wire buffer_auto_in_d_bits_source;
	wire buffer_auto_in_d_bits_sink;
	wire buffer_auto_in_d_bits_denied;
	wire [31:0] buffer_auto_in_d_bits_data;
	wire buffer_auto_in_d_bits_corrupt;
	wire buffer_auto_out_a_ready;
	wire buffer_auto_out_a_valid;
	wire [2:0] buffer_auto_out_a_bits_opcode;
	wire [2:0] buffer_auto_out_a_bits_param;
	wire [3:0] buffer_auto_out_a_bits_size;
	wire buffer_auto_out_a_bits_source;
	wire [31:0] buffer_auto_out_a_bits_address;
	wire [3:0] buffer_auto_out_a_bits_mask;
	wire [31:0] buffer_auto_out_a_bits_data;
	wire buffer_auto_out_a_bits_corrupt;
	wire buffer_auto_out_d_ready;
	wire buffer_auto_out_d_valid;
	wire [2:0] buffer_auto_out_d_bits_opcode;
	wire [1:0] buffer_auto_out_d_bits_param;
	wire [3:0] buffer_auto_out_d_bits_size;
	wire buffer_auto_out_d_bits_sink;
	wire buffer_auto_out_d_bits_denied;
	wire [31:0] buffer_auto_out_d_bits_data;
	wire buffer_auto_out_d_bits_corrupt;
	TLBuffer_5 buffer(
		.clock(buffer_clock),
		.reset(buffer_reset),
		.auto_in_a_ready(buffer_auto_in_a_ready),
		.auto_in_a_valid(buffer_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_auto_in_d_ready),
		.auto_in_d_valid(buffer_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_auto_out_a_ready),
		.auto_out_a_valid(buffer_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_auto_out_d_ready),
		.auto_out_d_valid(buffer_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(buffer_auto_out_d_bits_param),
		.auto_out_d_bits_size(buffer_auto_out_d_bits_size),
		.auto_out_d_bits_sink(buffer_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
		.auto_out_d_bits_data(buffer_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt)
	);
	assign auto_buffer_in_a_ready = buffer_auto_in_a_ready;
	assign auto_buffer_in_d_valid = buffer_auto_in_d_valid;
	assign auto_buffer_in_d_bits_opcode = buffer_auto_in_d_bits_opcode;
	assign auto_buffer_in_d_bits_param = buffer_auto_in_d_bits_param;
	assign auto_buffer_in_d_bits_size = buffer_auto_in_d_bits_size;
	assign auto_buffer_in_d_bits_source = buffer_auto_in_d_bits_source;
	assign auto_buffer_in_d_bits_sink = buffer_auto_in_d_bits_sink;
	assign auto_buffer_in_d_bits_denied = buffer_auto_in_d_bits_denied;
	assign auto_buffer_in_d_bits_data = buffer_auto_in_d_bits_data;
	assign auto_buffer_in_d_bits_corrupt = buffer_auto_in_d_bits_corrupt;
	assign auto_tl_out_a_valid = buffer_auto_out_a_valid;
	assign auto_tl_out_a_bits_opcode = buffer_auto_out_a_bits_opcode;
	assign auto_tl_out_a_bits_param = buffer_auto_out_a_bits_param;
	assign auto_tl_out_a_bits_size = buffer_auto_out_a_bits_size;
	assign auto_tl_out_a_bits_source = buffer_auto_out_a_bits_source;
	assign auto_tl_out_a_bits_address = buffer_auto_out_a_bits_address;
	assign auto_tl_out_a_bits_mask = buffer_auto_out_a_bits_mask;
	assign auto_tl_out_a_bits_data = buffer_auto_out_a_bits_data;
	assign auto_tl_out_a_bits_corrupt = buffer_auto_out_a_bits_corrupt;
	assign auto_tl_out_d_ready = buffer_auto_out_d_ready;
	assign buffer_clock = clock;
	assign buffer_reset = reset;
	assign buffer_auto_in_a_valid = auto_buffer_in_a_valid;
	assign buffer_auto_in_a_bits_opcode = auto_buffer_in_a_bits_opcode;
	assign buffer_auto_in_a_bits_param = auto_buffer_in_a_bits_param;
	assign buffer_auto_in_a_bits_size = auto_buffer_in_a_bits_size;
	assign buffer_auto_in_a_bits_source = auto_buffer_in_a_bits_source;
	assign buffer_auto_in_a_bits_address = auto_buffer_in_a_bits_address;
	assign buffer_auto_in_a_bits_mask = auto_buffer_in_a_bits_mask;
	assign buffer_auto_in_a_bits_data = auto_buffer_in_a_bits_data;
	assign buffer_auto_in_a_bits_corrupt = auto_buffer_in_a_bits_corrupt;
	assign buffer_auto_in_d_ready = auto_buffer_in_d_ready;
	assign buffer_auto_out_a_ready = auto_tl_out_a_ready;
	assign buffer_auto_out_d_valid = auto_tl_out_d_valid;
	assign buffer_auto_out_d_bits_opcode = auto_tl_out_d_bits_opcode;
	assign buffer_auto_out_d_bits_param = auto_tl_out_d_bits_param;
	assign buffer_auto_out_d_bits_size = auto_tl_out_d_bits_size;
	assign buffer_auto_out_d_bits_sink = auto_tl_out_d_bits_sink;
	assign buffer_auto_out_d_bits_denied = auto_tl_out_d_bits_denied;
	assign buffer_auto_out_d_bits_data = auto_tl_out_d_bits_data;
	assign buffer_auto_out_d_bits_corrupt = auto_tl_out_d_bits_corrupt;
endmodule
module FrontBus (
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_ready,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_valid,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_opcode,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_param,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_size,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_source,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_address,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_mask,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_data,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_corrupt,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_ready,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_valid,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_opcode,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_param,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_size,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_source,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_sink,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_denied,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_data,
	auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_corrupt,
	auto_fixedClockNode_out_clock,
	auto_fixedClockNode_out_reset,
	auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock,
	auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset,
	auto_bus_xing_out_a_ready,
	auto_bus_xing_out_a_valid,
	auto_bus_xing_out_a_bits_opcode,
	auto_bus_xing_out_a_bits_param,
	auto_bus_xing_out_a_bits_size,
	auto_bus_xing_out_a_bits_source,
	auto_bus_xing_out_a_bits_address,
	auto_bus_xing_out_a_bits_mask,
	auto_bus_xing_out_a_bits_data,
	auto_bus_xing_out_a_bits_corrupt,
	auto_bus_xing_out_d_ready,
	auto_bus_xing_out_d_valid,
	auto_bus_xing_out_d_bits_opcode,
	auto_bus_xing_out_d_bits_param,
	auto_bus_xing_out_d_bits_size,
	auto_bus_xing_out_d_bits_sink,
	auto_bus_xing_out_d_bits_denied,
	auto_bus_xing_out_d_bits_data,
	auto_bus_xing_out_d_bits_corrupt
);
	output wire auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_ready;
	input auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_valid;
	input [2:0] auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_opcode;
	input [2:0] auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_param;
	input [3:0] auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_size;
	input auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_source;
	input [31:0] auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_address;
	input [3:0] auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_mask;
	input [31:0] auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_data;
	input auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_corrupt;
	input auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_ready;
	output wire auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_valid;
	output wire [2:0] auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_opcode;
	output wire [1:0] auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_param;
	output wire [3:0] auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_size;
	output wire auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_source;
	output wire auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_sink;
	output wire auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_denied;
	output wire [31:0] auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_data;
	output wire auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_corrupt;
	output wire auto_fixedClockNode_out_clock;
	output wire auto_fixedClockNode_out_reset;
	input auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock;
	input auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset;
	input auto_bus_xing_out_a_ready;
	output wire auto_bus_xing_out_a_valid;
	output wire [2:0] auto_bus_xing_out_a_bits_opcode;
	output wire [2:0] auto_bus_xing_out_a_bits_param;
	output wire [3:0] auto_bus_xing_out_a_bits_size;
	output wire auto_bus_xing_out_a_bits_source;
	output wire [31:0] auto_bus_xing_out_a_bits_address;
	output wire [3:0] auto_bus_xing_out_a_bits_mask;
	output wire [31:0] auto_bus_xing_out_a_bits_data;
	output wire auto_bus_xing_out_a_bits_corrupt;
	output wire auto_bus_xing_out_d_ready;
	input auto_bus_xing_out_d_valid;
	input [2:0] auto_bus_xing_out_d_bits_opcode;
	input [1:0] auto_bus_xing_out_d_bits_param;
	input [3:0] auto_bus_xing_out_d_bits_size;
	input auto_bus_xing_out_d_bits_sink;
	input auto_bus_xing_out_d_bits_denied;
	input [31:0] auto_bus_xing_out_d_bits_data;
	input auto_bus_xing_out_d_bits_corrupt;
	wire subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_clock;
	wire subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_reset;
	wire subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_clock;
	wire subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_reset;
	wire clockGroup_auto_in_member_subsystem_fbus_0_clock;
	wire clockGroup_auto_in_member_subsystem_fbus_0_reset;
	wire clockGroup_auto_out_clock;
	wire clockGroup_auto_out_reset;
	wire fixedClockNode_auto_in_clock;
	wire fixedClockNode_auto_in_reset;
	wire fixedClockNode_auto_out_1_clock;
	wire fixedClockNode_auto_out_1_reset;
	wire fixedClockNode_auto_out_0_clock;
	wire fixedClockNode_auto_out_0_reset;
	wire subsystem_fbus_xbar_auto_in_a_ready;
	wire subsystem_fbus_xbar_auto_in_a_valid;
	wire [2:0] subsystem_fbus_xbar_auto_in_a_bits_opcode;
	wire [2:0] subsystem_fbus_xbar_auto_in_a_bits_param;
	wire [3:0] subsystem_fbus_xbar_auto_in_a_bits_size;
	wire subsystem_fbus_xbar_auto_in_a_bits_source;
	wire [31:0] subsystem_fbus_xbar_auto_in_a_bits_address;
	wire [3:0] subsystem_fbus_xbar_auto_in_a_bits_mask;
	wire [31:0] subsystem_fbus_xbar_auto_in_a_bits_data;
	wire subsystem_fbus_xbar_auto_in_a_bits_corrupt;
	wire subsystem_fbus_xbar_auto_in_d_ready;
	wire subsystem_fbus_xbar_auto_in_d_valid;
	wire [2:0] subsystem_fbus_xbar_auto_in_d_bits_opcode;
	wire [1:0] subsystem_fbus_xbar_auto_in_d_bits_param;
	wire [3:0] subsystem_fbus_xbar_auto_in_d_bits_size;
	wire subsystem_fbus_xbar_auto_in_d_bits_sink;
	wire subsystem_fbus_xbar_auto_in_d_bits_denied;
	wire [31:0] subsystem_fbus_xbar_auto_in_d_bits_data;
	wire subsystem_fbus_xbar_auto_in_d_bits_corrupt;
	wire subsystem_fbus_xbar_auto_out_a_ready;
	wire subsystem_fbus_xbar_auto_out_a_valid;
	wire [2:0] subsystem_fbus_xbar_auto_out_a_bits_opcode;
	wire [2:0] subsystem_fbus_xbar_auto_out_a_bits_param;
	wire [3:0] subsystem_fbus_xbar_auto_out_a_bits_size;
	wire subsystem_fbus_xbar_auto_out_a_bits_source;
	wire [31:0] subsystem_fbus_xbar_auto_out_a_bits_address;
	wire [3:0] subsystem_fbus_xbar_auto_out_a_bits_mask;
	wire [31:0] subsystem_fbus_xbar_auto_out_a_bits_data;
	wire subsystem_fbus_xbar_auto_out_a_bits_corrupt;
	wire subsystem_fbus_xbar_auto_out_d_ready;
	wire subsystem_fbus_xbar_auto_out_d_valid;
	wire [2:0] subsystem_fbus_xbar_auto_out_d_bits_opcode;
	wire [1:0] subsystem_fbus_xbar_auto_out_d_bits_param;
	wire [3:0] subsystem_fbus_xbar_auto_out_d_bits_size;
	wire subsystem_fbus_xbar_auto_out_d_bits_sink;
	wire subsystem_fbus_xbar_auto_out_d_bits_denied;
	wire [31:0] subsystem_fbus_xbar_auto_out_d_bits_data;
	wire subsystem_fbus_xbar_auto_out_d_bits_corrupt;
	wire buffer_clock;
	wire buffer_reset;
	wire buffer_auto_in_a_ready;
	wire buffer_auto_in_a_valid;
	wire [2:0] buffer_auto_in_a_bits_opcode;
	wire [2:0] buffer_auto_in_a_bits_param;
	wire [3:0] buffer_auto_in_a_bits_size;
	wire buffer_auto_in_a_bits_source;
	wire [31:0] buffer_auto_in_a_bits_address;
	wire [3:0] buffer_auto_in_a_bits_mask;
	wire [31:0] buffer_auto_in_a_bits_data;
	wire buffer_auto_in_a_bits_corrupt;
	wire buffer_auto_in_d_ready;
	wire buffer_auto_in_d_valid;
	wire [2:0] buffer_auto_in_d_bits_opcode;
	wire [1:0] buffer_auto_in_d_bits_param;
	wire [3:0] buffer_auto_in_d_bits_size;
	wire buffer_auto_in_d_bits_sink;
	wire buffer_auto_in_d_bits_denied;
	wire [31:0] buffer_auto_in_d_bits_data;
	wire buffer_auto_in_d_bits_corrupt;
	wire buffer_auto_out_a_ready;
	wire buffer_auto_out_a_valid;
	wire [2:0] buffer_auto_out_a_bits_opcode;
	wire [2:0] buffer_auto_out_a_bits_param;
	wire [3:0] buffer_auto_out_a_bits_size;
	wire buffer_auto_out_a_bits_source;
	wire [31:0] buffer_auto_out_a_bits_address;
	wire [3:0] buffer_auto_out_a_bits_mask;
	wire [31:0] buffer_auto_out_a_bits_data;
	wire buffer_auto_out_a_bits_corrupt;
	wire buffer_auto_out_d_ready;
	wire buffer_auto_out_d_valid;
	wire [2:0] buffer_auto_out_d_bits_opcode;
	wire [1:0] buffer_auto_out_d_bits_param;
	wire [3:0] buffer_auto_out_d_bits_size;
	wire buffer_auto_out_d_bits_sink;
	wire buffer_auto_out_d_bits_denied;
	wire [31:0] buffer_auto_out_d_bits_data;
	wire buffer_auto_out_d_bits_corrupt;
	wire coupler_from_port_named_serial_tl_ctrl_clock;
	wire coupler_from_port_named_serial_tl_ctrl_reset;
	wire coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_ready;
	wire coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_valid;
	wire [2:0] coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_opcode;
	wire [2:0] coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_param;
	wire [3:0] coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_size;
	wire coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_source;
	wire [31:0] coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_address;
	wire [3:0] coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_mask;
	wire [31:0] coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_data;
	wire coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_corrupt;
	wire coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_ready;
	wire coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_valid;
	wire [2:0] coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_opcode;
	wire [1:0] coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_param;
	wire [3:0] coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_size;
	wire coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_source;
	wire coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_sink;
	wire coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_denied;
	wire [31:0] coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_data;
	wire coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_corrupt;
	wire coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_ready;
	wire coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_valid;
	wire [2:0] coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_opcode;
	wire [2:0] coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_param;
	wire [3:0] coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_size;
	wire coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_source;
	wire [31:0] coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_address;
	wire [3:0] coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_mask;
	wire [31:0] coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_data;
	wire coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_corrupt;
	wire coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_ready;
	wire coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_valid;
	wire [2:0] coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_opcode;
	wire [1:0] coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_param;
	wire [3:0] coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_size;
	wire coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_sink;
	wire coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_denied;
	wire [31:0] coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_data;
	wire coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_corrupt;
	ClockGroupAggregator_2 subsystem_fbus_clock_groups(
		.auto_in_member_subsystem_fbus_0_clock(subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_clock),
		.auto_in_member_subsystem_fbus_0_reset(subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_reset),
		.auto_out_member_subsystem_fbus_0_clock(subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_clock),
		.auto_out_member_subsystem_fbus_0_reset(subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_reset)
	);
	ClockGroup_2 clockGroup(
		.auto_in_member_subsystem_fbus_0_clock(clockGroup_auto_in_member_subsystem_fbus_0_clock),
		.auto_in_member_subsystem_fbus_0_reset(clockGroup_auto_in_member_subsystem_fbus_0_reset),
		.auto_out_clock(clockGroup_auto_out_clock),
		.auto_out_reset(clockGroup_auto_out_reset)
	);
	FixedClockBroadcast_1 fixedClockNode(
		.auto_in_clock(fixedClockNode_auto_in_clock),
		.auto_in_reset(fixedClockNode_auto_in_reset),
		.auto_out_1_clock(fixedClockNode_auto_out_1_clock),
		.auto_out_1_reset(fixedClockNode_auto_out_1_reset),
		.auto_out_0_clock(fixedClockNode_auto_out_0_clock),
		.auto_out_0_reset(fixedClockNode_auto_out_0_reset)
	);
	TLXbar_3 subsystem_fbus_xbar(
		.auto_in_a_ready(subsystem_fbus_xbar_auto_in_a_ready),
		.auto_in_a_valid(subsystem_fbus_xbar_auto_in_a_valid),
		.auto_in_a_bits_opcode(subsystem_fbus_xbar_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(subsystem_fbus_xbar_auto_in_a_bits_param),
		.auto_in_a_bits_size(subsystem_fbus_xbar_auto_in_a_bits_size),
		.auto_in_a_bits_source(subsystem_fbus_xbar_auto_in_a_bits_source),
		.auto_in_a_bits_address(subsystem_fbus_xbar_auto_in_a_bits_address),
		.auto_in_a_bits_mask(subsystem_fbus_xbar_auto_in_a_bits_mask),
		.auto_in_a_bits_data(subsystem_fbus_xbar_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(subsystem_fbus_xbar_auto_in_a_bits_corrupt),
		.auto_in_d_ready(subsystem_fbus_xbar_auto_in_d_ready),
		.auto_in_d_valid(subsystem_fbus_xbar_auto_in_d_valid),
		.auto_in_d_bits_opcode(subsystem_fbus_xbar_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(subsystem_fbus_xbar_auto_in_d_bits_param),
		.auto_in_d_bits_size(subsystem_fbus_xbar_auto_in_d_bits_size),
		.auto_in_d_bits_sink(subsystem_fbus_xbar_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(subsystem_fbus_xbar_auto_in_d_bits_denied),
		.auto_in_d_bits_data(subsystem_fbus_xbar_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(subsystem_fbus_xbar_auto_in_d_bits_corrupt),
		.auto_out_a_ready(subsystem_fbus_xbar_auto_out_a_ready),
		.auto_out_a_valid(subsystem_fbus_xbar_auto_out_a_valid),
		.auto_out_a_bits_opcode(subsystem_fbus_xbar_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(subsystem_fbus_xbar_auto_out_a_bits_param),
		.auto_out_a_bits_size(subsystem_fbus_xbar_auto_out_a_bits_size),
		.auto_out_a_bits_source(subsystem_fbus_xbar_auto_out_a_bits_source),
		.auto_out_a_bits_address(subsystem_fbus_xbar_auto_out_a_bits_address),
		.auto_out_a_bits_mask(subsystem_fbus_xbar_auto_out_a_bits_mask),
		.auto_out_a_bits_data(subsystem_fbus_xbar_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(subsystem_fbus_xbar_auto_out_a_bits_corrupt),
		.auto_out_d_ready(subsystem_fbus_xbar_auto_out_d_ready),
		.auto_out_d_valid(subsystem_fbus_xbar_auto_out_d_valid),
		.auto_out_d_bits_opcode(subsystem_fbus_xbar_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(subsystem_fbus_xbar_auto_out_d_bits_param),
		.auto_out_d_bits_size(subsystem_fbus_xbar_auto_out_d_bits_size),
		.auto_out_d_bits_sink(subsystem_fbus_xbar_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(subsystem_fbus_xbar_auto_out_d_bits_denied),
		.auto_out_d_bits_data(subsystem_fbus_xbar_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(subsystem_fbus_xbar_auto_out_d_bits_corrupt)
	);
	TLBuffer_4 buffer(
		.clock(buffer_clock),
		.reset(buffer_reset),
		.auto_in_a_ready(buffer_auto_in_a_ready),
		.auto_in_a_valid(buffer_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_auto_in_d_ready),
		.auto_in_d_valid(buffer_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_auto_in_d_bits_size),
		.auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_auto_out_a_ready),
		.auto_out_a_valid(buffer_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_auto_out_d_ready),
		.auto_out_d_valid(buffer_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(buffer_auto_out_d_bits_param),
		.auto_out_d_bits_size(buffer_auto_out_d_bits_size),
		.auto_out_d_bits_sink(buffer_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
		.auto_out_d_bits_data(buffer_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt)
	);
	TLInterconnectCoupler_8 coupler_from_port_named_serial_tl_ctrl(
		.clock(coupler_from_port_named_serial_tl_ctrl_clock),
		.reset(coupler_from_port_named_serial_tl_ctrl_reset),
		.auto_buffer_in_a_ready(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_ready),
		.auto_buffer_in_a_valid(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_valid),
		.auto_buffer_in_a_bits_opcode(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_opcode),
		.auto_buffer_in_a_bits_param(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_param),
		.auto_buffer_in_a_bits_size(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_size),
		.auto_buffer_in_a_bits_source(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_source),
		.auto_buffer_in_a_bits_address(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_address),
		.auto_buffer_in_a_bits_mask(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_mask),
		.auto_buffer_in_a_bits_data(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_data),
		.auto_buffer_in_a_bits_corrupt(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_corrupt),
		.auto_buffer_in_d_ready(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_ready),
		.auto_buffer_in_d_valid(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_valid),
		.auto_buffer_in_d_bits_opcode(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_opcode),
		.auto_buffer_in_d_bits_param(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_param),
		.auto_buffer_in_d_bits_size(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_size),
		.auto_buffer_in_d_bits_source(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_source),
		.auto_buffer_in_d_bits_sink(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_sink),
		.auto_buffer_in_d_bits_denied(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_denied),
		.auto_buffer_in_d_bits_data(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_data),
		.auto_buffer_in_d_bits_corrupt(coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_corrupt),
		.auto_tl_out_a_ready(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_ready),
		.auto_tl_out_a_valid(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_valid),
		.auto_tl_out_a_bits_opcode(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_opcode),
		.auto_tl_out_a_bits_param(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_param),
		.auto_tl_out_a_bits_size(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_size),
		.auto_tl_out_a_bits_source(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_source),
		.auto_tl_out_a_bits_address(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_address),
		.auto_tl_out_a_bits_mask(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_mask),
		.auto_tl_out_a_bits_data(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_data),
		.auto_tl_out_a_bits_corrupt(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_corrupt),
		.auto_tl_out_d_ready(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_ready),
		.auto_tl_out_d_valid(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_valid),
		.auto_tl_out_d_bits_opcode(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_opcode),
		.auto_tl_out_d_bits_param(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_param),
		.auto_tl_out_d_bits_size(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_size),
		.auto_tl_out_d_bits_sink(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_sink),
		.auto_tl_out_d_bits_denied(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_denied),
		.auto_tl_out_d_bits_data(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_data),
		.auto_tl_out_d_bits_corrupt(coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_corrupt)
	);
	assign auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_ready = coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_ready;
	assign auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_valid = coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_valid;
	assign auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_opcode = coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_opcode;
	assign auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_param = coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_param;
	assign auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_size = coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_size;
	assign auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_source = coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_source;
	assign auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_sink = coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_sink;
	assign auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_denied = coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_denied;
	assign auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_data = coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_data;
	assign auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_corrupt = coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_bits_corrupt;
	assign auto_fixedClockNode_out_clock = fixedClockNode_auto_out_1_clock;
	assign auto_fixedClockNode_out_reset = fixedClockNode_auto_out_1_reset;
	assign auto_bus_xing_out_a_valid = buffer_auto_out_a_valid;
	assign auto_bus_xing_out_a_bits_opcode = buffer_auto_out_a_bits_opcode;
	assign auto_bus_xing_out_a_bits_param = buffer_auto_out_a_bits_param;
	assign auto_bus_xing_out_a_bits_size = buffer_auto_out_a_bits_size;
	assign auto_bus_xing_out_a_bits_source = buffer_auto_out_a_bits_source;
	assign auto_bus_xing_out_a_bits_address = buffer_auto_out_a_bits_address;
	assign auto_bus_xing_out_a_bits_mask = buffer_auto_out_a_bits_mask;
	assign auto_bus_xing_out_a_bits_data = buffer_auto_out_a_bits_data;
	assign auto_bus_xing_out_a_bits_corrupt = buffer_auto_out_a_bits_corrupt;
	assign auto_bus_xing_out_d_ready = buffer_auto_out_d_ready;
	assign subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_clock = auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock;
	assign subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_reset = auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset;
	assign clockGroup_auto_in_member_subsystem_fbus_0_clock = subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_clock;
	assign clockGroup_auto_in_member_subsystem_fbus_0_reset = subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_reset;
	assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock;
	assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset;
	assign subsystem_fbus_xbar_auto_in_a_valid = coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_valid;
	assign subsystem_fbus_xbar_auto_in_a_bits_opcode = coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_opcode;
	assign subsystem_fbus_xbar_auto_in_a_bits_param = coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_param;
	assign subsystem_fbus_xbar_auto_in_a_bits_size = coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_size;
	assign subsystem_fbus_xbar_auto_in_a_bits_source = coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_source;
	assign subsystem_fbus_xbar_auto_in_a_bits_address = coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_address;
	assign subsystem_fbus_xbar_auto_in_a_bits_mask = coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_mask;
	assign subsystem_fbus_xbar_auto_in_a_bits_data = coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_data;
	assign subsystem_fbus_xbar_auto_in_a_bits_corrupt = coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_bits_corrupt;
	assign subsystem_fbus_xbar_auto_in_d_ready = coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_ready;
	assign subsystem_fbus_xbar_auto_out_a_ready = buffer_auto_in_a_ready;
	assign subsystem_fbus_xbar_auto_out_d_valid = buffer_auto_in_d_valid;
	assign subsystem_fbus_xbar_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode;
	assign subsystem_fbus_xbar_auto_out_d_bits_param = buffer_auto_in_d_bits_param;
	assign subsystem_fbus_xbar_auto_out_d_bits_size = buffer_auto_in_d_bits_size;
	assign subsystem_fbus_xbar_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink;
	assign subsystem_fbus_xbar_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied;
	assign subsystem_fbus_xbar_auto_out_d_bits_data = buffer_auto_in_d_bits_data;
	assign subsystem_fbus_xbar_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt;
	assign buffer_clock = fixedClockNode_auto_out_0_clock;
	assign buffer_reset = fixedClockNode_auto_out_0_reset;
	assign buffer_auto_in_a_valid = subsystem_fbus_xbar_auto_out_a_valid;
	assign buffer_auto_in_a_bits_opcode = subsystem_fbus_xbar_auto_out_a_bits_opcode;
	assign buffer_auto_in_a_bits_param = subsystem_fbus_xbar_auto_out_a_bits_param;
	assign buffer_auto_in_a_bits_size = subsystem_fbus_xbar_auto_out_a_bits_size;
	assign buffer_auto_in_a_bits_source = subsystem_fbus_xbar_auto_out_a_bits_source;
	assign buffer_auto_in_a_bits_address = subsystem_fbus_xbar_auto_out_a_bits_address;
	assign buffer_auto_in_a_bits_mask = subsystem_fbus_xbar_auto_out_a_bits_mask;
	assign buffer_auto_in_a_bits_data = subsystem_fbus_xbar_auto_out_a_bits_data;
	assign buffer_auto_in_a_bits_corrupt = subsystem_fbus_xbar_auto_out_a_bits_corrupt;
	assign buffer_auto_in_d_ready = subsystem_fbus_xbar_auto_out_d_ready;
	assign buffer_auto_out_a_ready = auto_bus_xing_out_a_ready;
	assign buffer_auto_out_d_valid = auto_bus_xing_out_d_valid;
	assign buffer_auto_out_d_bits_opcode = auto_bus_xing_out_d_bits_opcode;
	assign buffer_auto_out_d_bits_param = auto_bus_xing_out_d_bits_param;
	assign buffer_auto_out_d_bits_size = auto_bus_xing_out_d_bits_size;
	assign buffer_auto_out_d_bits_sink = auto_bus_xing_out_d_bits_sink;
	assign buffer_auto_out_d_bits_denied = auto_bus_xing_out_d_bits_denied;
	assign buffer_auto_out_d_bits_data = auto_bus_xing_out_d_bits_data;
	assign buffer_auto_out_d_bits_corrupt = auto_bus_xing_out_d_bits_corrupt;
	assign coupler_from_port_named_serial_tl_ctrl_clock = fixedClockNode_auto_out_0_clock;
	assign coupler_from_port_named_serial_tl_ctrl_reset = fixedClockNode_auto_out_0_reset;
	assign coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_valid = auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_valid;
	assign coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_opcode = auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_opcode;
	assign coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_param = auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_param;
	assign coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_size = auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_size;
	assign coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_source = auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_source;
	assign coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_address = auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_address;
	assign coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_mask = auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_mask;
	assign coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_data = auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_data;
	assign coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_a_bits_corrupt = auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_corrupt;
	assign coupler_from_port_named_serial_tl_ctrl_auto_buffer_in_d_ready = auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_ready;
	assign coupler_from_port_named_serial_tl_ctrl_auto_tl_out_a_ready = subsystem_fbus_xbar_auto_in_a_ready;
	assign coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_valid = subsystem_fbus_xbar_auto_in_d_valid;
	assign coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_opcode = subsystem_fbus_xbar_auto_in_d_bits_opcode;
	assign coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_param = subsystem_fbus_xbar_auto_in_d_bits_param;
	assign coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_size = subsystem_fbus_xbar_auto_in_d_bits_size;
	assign coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_sink = subsystem_fbus_xbar_auto_in_d_bits_sink;
	assign coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_denied = subsystem_fbus_xbar_auto_in_d_bits_denied;
	assign coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_data = subsystem_fbus_xbar_auto_in_d_bits_data;
	assign coupler_from_port_named_serial_tl_ctrl_auto_tl_out_d_bits_corrupt = subsystem_fbus_xbar_auto_in_d_bits_corrupt;
endmodule
module ClockGroupAggregator_3 (
	auto_in_member_subsystem_cbus_0_clock,
	auto_in_member_subsystem_cbus_0_reset,
	auto_out_member_subsystem_cbus_0_clock,
	auto_out_member_subsystem_cbus_0_reset
);
	input auto_in_member_subsystem_cbus_0_clock;
	input auto_in_member_subsystem_cbus_0_reset;
	output wire auto_out_member_subsystem_cbus_0_clock;
	output wire auto_out_member_subsystem_cbus_0_reset;
	assign auto_out_member_subsystem_cbus_0_clock = auto_in_member_subsystem_cbus_0_clock;
	assign auto_out_member_subsystem_cbus_0_reset = auto_in_member_subsystem_cbus_0_reset;
endmodule
module ClockGroup_3 (
	auto_in_member_subsystem_cbus_0_clock,
	auto_in_member_subsystem_cbus_0_reset,
	auto_out_clock,
	auto_out_reset
);
	input auto_in_member_subsystem_cbus_0_clock;
	input auto_in_member_subsystem_cbus_0_reset;
	output wire auto_out_clock;
	output wire auto_out_reset;
	assign auto_out_clock = auto_in_member_subsystem_cbus_0_clock;
	assign auto_out_reset = auto_in_member_subsystem_cbus_0_reset;
endmodule
module FixedClockBroadcast_3 (
	auto_in_clock,
	auto_in_reset,
	auto_out_5_clock,
	auto_out_5_reset,
	auto_out_4_clock,
	auto_out_4_reset,
	auto_out_3_clock,
	auto_out_3_reset,
	auto_out_1_clock,
	auto_out_1_reset,
	auto_out_0_clock,
	auto_out_0_reset
);
	input auto_in_clock;
	input auto_in_reset;
	output wire auto_out_5_clock;
	output wire auto_out_5_reset;
	output wire auto_out_4_clock;
	output wire auto_out_4_reset;
	output wire auto_out_3_clock;
	output wire auto_out_3_reset;
	output wire auto_out_1_clock;
	output wire auto_out_1_reset;
	output wire auto_out_0_clock;
	output wire auto_out_0_reset;
	assign auto_out_5_clock = auto_in_clock;
	assign auto_out_5_reset = auto_in_reset;
	assign auto_out_4_clock = auto_in_clock;
	assign auto_out_4_reset = auto_in_reset;
	assign auto_out_3_clock = auto_in_clock;
	assign auto_out_3_reset = auto_in_reset;
	assign auto_out_1_clock = auto_in_clock;
	assign auto_out_1_reset = auto_in_reset;
	assign auto_out_0_clock = auto_in_clock;
	assign auto_out_0_reset = auto_in_reset;
endmodule
module TLMonitor_15 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire _T_44 = io_in_a_bits_size <= 4'hc;
	wire _T_53 = _T_44 & source_ok;
	wire [32:0] _T_59 = $signed(_T_7) & -33'sh000005000;
	wire _T_60 = $signed(_T_59) == 33'sh000000000;
	wire [31:0] _T_61 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_62 = {1'b0, $signed(_T_61)};
	wire [32:0] _T_64 = $signed(_T_62) & -33'sh000001000;
	wire _T_65 = $signed(_T_64) == 33'sh000000000;
	wire [31:0] _T_66 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_67 = {1'b0, $signed(_T_66)};
	wire [32:0] _T_69 = $signed(_T_67) & -33'sh000010000;
	wire _T_70 = $signed(_T_69) == 33'sh000000000;
	wire [31:0] _T_71 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_72 = {1'b0, $signed(_T_71)};
	wire [32:0] _T_74 = $signed(_T_72) & -33'sh000010000;
	wire _T_75 = $signed(_T_74) == 33'sh000000000;
	wire [31:0] _T_76 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_77 = {1'b0, $signed(_T_76)};
	wire [32:0] _T_79 = $signed(_T_77) & -33'sh000011000;
	wire _T_80 = $signed(_T_79) == 33'sh000000000;
	wire [31:0] _T_81 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_82 = {1'b0, $signed(_T_81)};
	wire [32:0] _T_84 = $signed(_T_82) & -33'sh000010000;
	wire _T_85 = $signed(_T_84) == 33'sh000000000;
	wire [31:0] _T_86 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_87 = {1'b0, $signed(_T_86)};
	wire [32:0] _T_89 = $signed(_T_87) & -33'sh004000000;
	wire _T_90 = $signed(_T_89) == 33'sh000000000;
	wire [31:0] _T_91 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_92 = {1'b0, $signed(_T_91)};
	wire [32:0] _T_94 = $signed(_T_92) & -33'sh000001000;
	wire _T_95 = $signed(_T_94) == 33'sh000000000;
	wire [31:0] _T_96 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_97 = {1'b0, $signed(_T_96)};
	wire [32:0] _T_99 = $signed(_T_97) & -33'sh000001000;
	wire _T_100 = $signed(_T_99) == 33'sh000000000;
	wire [31:0] _T_101 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_102 = {1'b0, $signed(_T_101)};
	wire [32:0] _T_104 = $signed(_T_102) & -33'sh000004000;
	wire _T_105 = $signed(_T_104) == 33'sh000000000;
	wire _T_200 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_204 = ~io_in_a_bits_mask;
	wire _T_205 = _T_204 == 4'h0;
	wire _T_209 = ~io_in_a_bits_corrupt;
	wire _T_213 = io_in_a_bits_opcode == 3'h7;
	wire _T_375 = io_in_a_bits_param != 3'h0;
	wire _T_388 = io_in_a_bits_opcode == 3'h4;
	wire _T_413 = _T_44 & _T_65;
	wire _T_415 = io_in_a_bits_size <= 4'h6;
	wire _T_470 = (((((((_T_60 | _T_70) | _T_75) | _T_80) | _T_85) | _T_90) | _T_95) | _T_100) | _T_105;
	wire _T_471 = _T_415 & _T_470;
	wire _T_473 = _T_413 | _T_471;
	wire _T_483 = io_in_a_bits_param == 3'h0;
	wire _T_487 = io_in_a_bits_mask == mask;
	wire _T_495 = io_in_a_bits_opcode == 3'h0;
	wire _T_562 = (((((_T_60 | _T_80) | _T_85) | _T_90) | _T_95) | _T_100) | _T_105;
	wire _T_563 = _T_415 & _T_562;
	wire _T_578 = _T_413 | _T_563;
	wire _T_580 = _T_53 & _T_578;
	wire _T_598 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_697 = ~mask;
	wire [3:0] _T_698 = io_in_a_bits_mask & _T_697;
	wire _T_699 = _T_698 == 4'h0;
	wire _T_703 = io_in_a_bits_opcode == 3'h2;
	wire _T_717 = io_in_a_bits_size <= 4'h2;
	wire [31:0] _T_725 = io_in_a_bits_address ^ 32'h00004000;
	wire [32:0] _T_726 = {1'b0, $signed(_T_725)};
	wire [32:0] _T_728 = $signed(_T_726) & -33'sh000001000;
	wire _T_729 = $signed(_T_728) == 33'sh000000000;
	wire _T_742 = ((_T_65 | _T_729) | _T_95) | _T_100;
	wire _T_743 = _T_717 & _T_742;
	wire _T_781 = 4'h2 == io_in_a_bits_size;
	wire _T_788 = _T_781 & _T_105;
	wire _T_791 = _T_743 | _T_788;
	wire _T_792 = _T_53 & _T_791;
	wire _T_802 = io_in_a_bits_param <= 3'h4;
	wire _T_810 = io_in_a_bits_opcode == 3'h3;
	wire _T_909 = io_in_a_bits_param <= 3'h3;
	wire _T_917 = io_in_a_bits_opcode == 3'h5;
	wire _T_997 = _T_53 & _T_413;
	wire _T_1007 = io_in_a_bits_param <= 3'h1;
	wire _T_1019 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_1023 = io_in_d_bits_opcode == 3'h6;
	wire _T_1027 = io_in_d_bits_size >= 4'h2;
	wire _T_1031 = io_in_d_bits_param == 2'h0;
	wire _T_1035 = ~io_in_d_bits_corrupt;
	wire _T_1039 = ~io_in_d_bits_denied;
	wire _T_1043 = io_in_d_bits_opcode == 3'h4;
	wire _T_1054 = io_in_d_bits_param <= 2'h2;
	wire _T_1058 = io_in_d_bits_param != 2'h2;
	wire _T_1071 = io_in_d_bits_opcode == 3'h5;
	wire _T_1091 = _T_1039 | io_in_d_bits_corrupt;
	wire _T_1100 = io_in_d_bits_opcode == 3'h0;
	wire _T_1117 = io_in_d_bits_opcode == 3'h1;
	wire _T_1135 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg [2:0] source;
	reg [31:0] address;
	wire _T_1165 = io_in_a_valid & ~a_first;
	wire _T_1166 = io_in_a_bits_opcode == opcode;
	wire _T_1170 = io_in_a_bits_param == param;
	wire _T_1174 = io_in_a_bits_size == size;
	wire _T_1178 = io_in_a_bits_source == source;
	wire _T_1182 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_1189 = io_in_d_valid & ~d_first;
	wire _T_1190 = io_in_d_bits_opcode == opcode_1;
	wire _T_1194 = io_in_d_bits_param == param_1;
	wire _T_1198 = io_in_d_bits_size == size_1;
	wire _T_1202 = io_in_d_bits_source == source_1;
	wire _T_1206 = io_in_d_bits_sink == sink;
	wire _T_1210 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [39:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [5:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0};
	wire [39:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T;
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [39:0] _GEN_75 = {24'd0, _a_size_lookup_T_5};
	wire [39:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_75;
	wire [39:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[39:1]};
	wire _T_1216 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire _T_1219 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [4:0] _GEN_77 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_77};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [5:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [67:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [67:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire [4:0] _T_1221 = inflight >> io_in_a_bits_source;
	wire _T_1223 = ~_T_1221[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [67:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 68'h00000000000000000);
	wire _T_1227 = io_in_d_valid & d_first_1;
	wire _T_1229 = ~_T_1023;
	wire _T_1230 = (io_in_d_valid & d_first_1) & ~_T_1023;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [78:0] _GEN_4 = {63'd0, _a_size_lookup_T_5};
	wire [78:0] _d_sizes_clr_T_5 = _GEN_4 << _a_size_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_1229 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1229 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [78:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1229 ? _d_sizes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_1216 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_1240 = inflight >> io_in_d_bits_source;
	wire _T_1242 = _T_1240[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1247 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1248 = (io_in_d_bits_opcode == _GEN_32) | _T_1247;
	wire _T_1252 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1259 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1260 = (io_in_d_bits_opcode == _GEN_48) | _T_1259;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_79 = {4'd0, io_in_d_bits_size};
	wire _T_1264 = _GEN_79 == a_size_lookup;
	wire _T_1274 = (((_T_1227 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_1229;
	wire _T_1276 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [39:0] a_sizes_set = _GEN_20[39:0];
	wire [39:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [39:0] d_sizes_clr = _GEN_24[39:0];
	wire [39:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [39:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1285 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [39:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [39:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T;
	wire [39:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_75;
	wire [39:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[39:1]};
	wire _T_1311 = (io_in_d_valid & d_first_2) & _T_1023;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_1023 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_1023 ? _d_sizes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_1319 = inflight_1 >> io_in_d_bits_source;
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1329 = _GEN_79 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [39:0] d_sizes_clr_1 = _GEN_69[39:0];
	wire [39:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [39:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	reg [31:0] watchdog_1;
	wire _T_1349 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 40'h0000000000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 40'h0000000000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLFIFOFixer_2 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [31:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [3:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	TLMonitor_15 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_out_a_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid;
	assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_io_in_d_bits_param = auto_out_d_bits_param;
	assign monitor_io_in_d_bits_size = auto_out_d_bits_size;
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source;
	assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink;
	assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied;
	assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt;
endmodule
module TLMonitor_16 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input [1:0] io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input [1:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 2'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 2'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 2'h0;
	wire source_ok = (_source_ok_T | _source_ok_T_1) | _source_ok_T_2;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_33 = io_in_a_bits_opcode == 3'h6;
	wire _T_35 = io_in_a_bits_size <= 4'hc;
	wire _T_42 = _T_35 & source_ok;
	wire [32:0] _T_48 = $signed(_T_7) & -33'sh000005000;
	wire _T_49 = $signed(_T_48) == 33'sh000000000;
	wire [31:0] _T_50 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_51 = {1'b0, $signed(_T_50)};
	wire [32:0] _T_53 = $signed(_T_51) & -33'sh000001000;
	wire _T_54 = $signed(_T_53) == 33'sh000000000;
	wire [31:0] _T_55 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_56 = {1'b0, $signed(_T_55)};
	wire [32:0] _T_58 = $signed(_T_56) & -33'sh000010000;
	wire _T_59 = $signed(_T_58) == 33'sh000000000;
	wire [31:0] _T_60 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_61 = {1'b0, $signed(_T_60)};
	wire [32:0] _T_63 = $signed(_T_61) & -33'sh000010000;
	wire _T_64 = $signed(_T_63) == 33'sh000000000;
	wire [31:0] _T_65 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_66 = {1'b0, $signed(_T_65)};
	wire [32:0] _T_68 = $signed(_T_66) & -33'sh000011000;
	wire _T_69 = $signed(_T_68) == 33'sh000000000;
	wire [31:0] _T_70 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_71 = {1'b0, $signed(_T_70)};
	wire [32:0] _T_73 = $signed(_T_71) & -33'sh000010000;
	wire _T_74 = $signed(_T_73) == 33'sh000000000;
	wire [31:0] _T_75 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_76 = {1'b0, $signed(_T_75)};
	wire [32:0] _T_78 = $signed(_T_76) & -33'sh004000000;
	wire _T_79 = $signed(_T_78) == 33'sh000000000;
	wire [31:0] _T_80 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_81 = {1'b0, $signed(_T_80)};
	wire [32:0] _T_83 = $signed(_T_81) & -33'sh000001000;
	wire _T_84 = $signed(_T_83) == 33'sh000000000;
	wire [31:0] _T_85 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_86 = {1'b0, $signed(_T_85)};
	wire [32:0] _T_88 = $signed(_T_86) & -33'sh000001000;
	wire _T_89 = $signed(_T_88) == 33'sh000000000;
	wire [31:0] _T_90 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_91 = {1'b0, $signed(_T_90)};
	wire [32:0] _T_93 = $signed(_T_91) & -33'sh000004000;
	wire _T_94 = $signed(_T_93) == 33'sh000000000;
	wire _T_189 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_193 = ~io_in_a_bits_mask;
	wire _T_194 = _T_193 == 4'h0;
	wire _T_198 = ~io_in_a_bits_corrupt;
	wire _T_202 = io_in_a_bits_opcode == 3'h7;
	wire _T_362 = io_in_a_bits_param != 3'h0;
	wire _T_375 = io_in_a_bits_opcode == 3'h4;
	wire _T_398 = _T_35 & _T_54;
	wire _T_400 = io_in_a_bits_size <= 4'h6;
	wire _T_455 = (((((((_T_49 | _T_59) | _T_64) | _T_69) | _T_74) | _T_79) | _T_84) | _T_89) | _T_94;
	wire _T_456 = _T_400 & _T_455;
	wire _T_458 = _T_398 | _T_456;
	wire _T_468 = io_in_a_bits_param == 3'h0;
	wire _T_472 = io_in_a_bits_mask == mask;
	wire _T_480 = io_in_a_bits_opcode == 3'h0;
	wire _T_545 = (((((_T_49 | _T_69) | _T_74) | _T_79) | _T_84) | _T_89) | _T_94;
	wire _T_546 = _T_400 & _T_545;
	wire _T_561 = _T_398 | _T_546;
	wire _T_563 = _T_42 & _T_561;
	wire _T_581 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_678 = ~mask;
	wire [3:0] _T_679 = io_in_a_bits_mask & _T_678;
	wire _T_680 = _T_679 == 4'h0;
	wire _T_684 = io_in_a_bits_opcode == 3'h2;
	wire _T_696 = io_in_a_bits_size <= 4'h2;
	wire _T_745 = ((((((_T_49 | _T_54) | _T_69) | _T_74) | _T_79) | _T_84) | _T_89) | _T_94;
	wire _T_746 = _T_696 & _T_745;
	wire _T_762 = _T_42 & _T_746;
	wire _T_772 = io_in_a_bits_param <= 3'h4;
	wire _T_780 = io_in_a_bits_opcode == 3'h3;
	wire _T_868 = io_in_a_bits_param <= 3'h3;
	wire _T_876 = io_in_a_bits_opcode == 3'h5;
	wire _T_954 = _T_42 & _T_398;
	wire _T_964 = io_in_a_bits_param <= 3'h1;
	wire _T_976 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_4 = io_in_d_bits_source == 2'h2;
	wire _source_ok_T_5 = io_in_d_bits_source == 2'h1;
	wire _source_ok_T_6 = io_in_d_bits_source == 2'h0;
	wire source_ok_1 = (_source_ok_T_4 | _source_ok_T_5) | _source_ok_T_6;
	wire _T_980 = io_in_d_bits_opcode == 3'h6;
	wire _T_984 = io_in_d_bits_size >= 4'h2;
	wire _T_988 = io_in_d_bits_param == 2'h0;
	wire _T_992 = ~io_in_d_bits_corrupt;
	wire _T_996 = ~io_in_d_bits_denied;
	wire _T_1000 = io_in_d_bits_opcode == 3'h4;
	wire _T_1011 = io_in_d_bits_param <= 2'h2;
	wire _T_1015 = io_in_d_bits_param != 2'h2;
	wire _T_1028 = io_in_d_bits_opcode == 3'h5;
	wire _T_1048 = _T_996 | io_in_d_bits_corrupt;
	wire _T_1057 = io_in_d_bits_opcode == 3'h0;
	wire _T_1074 = io_in_d_bits_opcode == 3'h1;
	wire _T_1092 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg [1:0] source;
	reg [31:0] address;
	wire _T_1122 = io_in_a_valid & ~a_first;
	wire _T_1123 = io_in_a_bits_opcode == opcode;
	wire _T_1127 = io_in_a_bits_param == param;
	wire _T_1131 = io_in_a_bits_size == size;
	wire _T_1135 = io_in_a_bits_source == source;
	wire _T_1139 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg [1:0] source_1;
	reg sink;
	reg denied;
	wire _T_1146 = io_in_d_valid & ~d_first;
	wire _T_1147 = io_in_d_bits_opcode == opcode_1;
	wire _T_1151 = io_in_d_bits_param == param_1;
	wire _T_1155 = io_in_d_bits_size == size_1;
	wire _T_1159 = io_in_d_bits_source == source_1;
	wire _T_1163 = io_in_d_bits_sink == sink;
	wire _T_1167 = io_in_d_bits_denied == denied;
	reg [2:0] inflight;
	reg [11:0] inflight_opcodes;
	reg [23:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [3:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [4:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [11:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_1};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [4:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0};
	wire [23:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T;
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [23:0] _GEN_75 = {8'd0, _a_size_lookup_T_5};
	wire [23:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_75;
	wire [23:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[23:1]};
	wire _T_1173 = io_in_a_valid & a_first_1;
	wire [3:0] _a_set_wo_ready_T = 4'h1 << io_in_a_bits_source;
	wire [3:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 4'h0);
	wire _T_1176 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [3:0] _GEN_77 = {io_in_a_bits_source, 2'h0};
	wire [4:0] _a_opcodes_set_T = {1'd0, _GEN_77};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [34:0] _GEN_1 = {31'd0, a_opcodes_set_interm};
	wire [34:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [4:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [35:0] _GEN_2 = {31'd0, a_sizes_set_interm};
	wire [35:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire [2:0] _T_1178 = inflight >> io_in_a_bits_source;
	wire _T_1180 = ~_T_1178[0];
	wire [3:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 4'h0);
	wire [34:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 35'h000000000);
	wire [35:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 36'h000000000);
	wire _T_1184 = io_in_d_valid & d_first_1;
	wire _T_1186 = ~_T_980;
	wire _T_1187 = (io_in_d_valid & d_first_1) & ~_T_980;
	wire [3:0] _d_clr_wo_ready_T = 4'h1 << io_in_d_bits_source;
	wire [3:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_980 ? _d_clr_wo_ready_T : 4'h0);
	wire [46:0] _GEN_3 = {31'd0, _a_opcode_lookup_T_5};
	wire [46:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [46:0] _GEN_4 = {31'd0, _a_size_lookup_T_5};
	wire [46:0] _d_sizes_clr_T_5 = _GEN_4 << _a_size_lookup_T;
	wire [3:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_1186 ? _d_clr_wo_ready_T : 4'h0);
	wire [46:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1186 ? _d_opcodes_clr_T_5 : 47'h000000000000);
	wire [46:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1186 ? _d_sizes_clr_T_5 : 47'h000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_1173 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [2:0] _T_1197 = inflight >> io_in_d_bits_source;
	wire _T_1199 = _T_1197[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1204 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1205 = (io_in_d_bits_opcode == _GEN_32) | _T_1204;
	wire _T_1209 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1216 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1217 = (io_in_d_bits_opcode == _GEN_48) | _T_1216;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_79 = {4'd0, io_in_d_bits_size};
	wire _T_1221 = _GEN_79 == a_size_lookup;
	wire _T_1231 = (((_T_1184 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_1186;
	wire _T_1233 = ~io_in_d_ready | io_in_a_ready;
	wire [2:0] a_set_wo_ready = _GEN_15[2:0];
	wire [2:0] d_clr_wo_ready = _GEN_21[2:0];
	wire _T_1240 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [2:0] a_set = _GEN_16[2:0];
	wire [2:0] _inflight_T = inflight | a_set;
	wire [2:0] d_clr = _GEN_22[2:0];
	wire [2:0] _inflight_T_1 = ~d_clr;
	wire [2:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [11:0] a_opcodes_set = _GEN_19[11:0];
	wire [11:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [11:0] d_opcodes_clr = _GEN_23[11:0];
	wire [11:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [11:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [23:0] a_sizes_set = _GEN_20[23:0];
	wire [23:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [23:0] d_sizes_clr = _GEN_24[23:0];
	wire [23:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [23:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1249 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [2:0] inflight_1;
	reg [23:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [23:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T;
	wire [23:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_75;
	wire [23:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[23:1]};
	wire _T_1275 = (io_in_d_valid & d_first_2) & _T_980;
	wire [3:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_980 ? _d_clr_wo_ready_T : 4'h0);
	wire [46:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_980 ? _d_sizes_clr_T_5 : 47'h000000000000);
	wire [2:0] _T_1283 = inflight_1 >> io_in_d_bits_source;
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1293 = _GEN_79 == c_size_lookup;
	wire [2:0] d_clr_1 = _GEN_67[2:0];
	wire [2:0] _inflight_T_4 = ~d_clr_1;
	wire [2:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [23:0] d_sizes_clr_1 = _GEN_69[23:0];
	wire [23:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [23:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	reg [31:0] watchdog_1;
	wire _T_1318 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 3'h0;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 12'h000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 24'h000000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 3'h0;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 24'h000000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLMonitor_17 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_address,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [31:0] io_in_a_bits_address;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire [31:0] _is_aligned_T = io_in_a_bits_address & 32'h00000003;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire [32:0] _T_26 = $signed(_T_7) & -33'sh000005000;
	wire _T_27 = $signed(_T_26) == 33'sh000000000;
	wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_29 = {1'b0, $signed(_T_28)};
	wire [32:0] _T_31 = $signed(_T_29) & -33'sh000001000;
	wire _T_32 = $signed(_T_31) == 33'sh000000000;
	wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_44 = {1'b0, $signed(_T_43)};
	wire [32:0] _T_46 = $signed(_T_44) & -33'sh000011000;
	wire _T_47 = $signed(_T_46) == 33'sh000000000;
	wire [31:0] _T_48 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_49 = {1'b0, $signed(_T_48)};
	wire [32:0] _T_51 = $signed(_T_49) & -33'sh000010000;
	wire _T_52 = $signed(_T_51) == 33'sh000000000;
	wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_54 = {1'b0, $signed(_T_53)};
	wire [32:0] _T_56 = $signed(_T_54) & -33'sh004000000;
	wire _T_57 = $signed(_T_56) == 33'sh000000000;
	wire [31:0] _T_58 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_59 = {1'b0, $signed(_T_58)};
	wire [32:0] _T_61 = $signed(_T_59) & -33'sh000001000;
	wire _T_62 = $signed(_T_61) == 33'sh000000000;
	wire [31:0] _T_63 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_64 = {1'b0, $signed(_T_63)};
	wire [32:0] _T_66 = $signed(_T_64) & -33'sh000001000;
	wire _T_67 = $signed(_T_66) == 33'sh000000000;
	wire [31:0] _T_68 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_69 = {1'b0, $signed(_T_68)};
	wire [32:0] _T_71 = $signed(_T_69) & -33'sh000004000;
	wire _T_72 = $signed(_T_71) == 33'sh000000000;
	wire _T_511 = (((((_T_27 | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_527 = _T_32 | _T_511;
	wire _T_926 = io_in_d_bits_opcode <= 3'h6;
	wire _T_930 = io_in_d_bits_opcode == 3'h6;
	wire _T_934 = io_in_d_bits_size >= 4'h2;
	wire _T_938 = io_in_d_bits_param == 2'h0;
	wire _T_942 = ~io_in_d_bits_corrupt;
	wire _T_946 = ~io_in_d_bits_denied;
	wire _T_950 = io_in_d_bits_opcode == 3'h4;
	wire _T_961 = io_in_d_bits_param <= 2'h2;
	wire _T_965 = io_in_d_bits_param != 2'h2;
	wire _T_978 = io_in_d_bits_opcode == 3'h5;
	wire _T_998 = _T_946 | io_in_d_bits_corrupt;
	wire _T_1007 = io_in_d_bits_opcode == 3'h0;
	wire _T_1024 = io_in_d_bits_opcode == 3'h1;
	wire _T_1042 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [31:0] address;
	wire _T_1072 = io_in_a_valid & ~a_first;
	wire _T_1089 = io_in_a_bits_address == address;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg sink;
	reg denied;
	wire _T_1096 = io_in_d_valid & ~d_first;
	wire _T_1097 = io_in_d_bits_opcode == opcode_1;
	wire _T_1101 = io_in_d_bits_param == param_1;
	wire _T_1105 = io_in_d_bits_size == size_1;
	wire _T_1113 = io_in_d_bits_sink == sink;
	wire _T_1117 = io_in_d_bits_denied == denied;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [7:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_71 = {12'd0, inflight_opcodes};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_71 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [15:0] _GEN_73 = {8'd0, inflight_sizes};
	wire [15:0] _a_size_lookup_T_6 = _GEN_73 & _a_size_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_1123 = io_in_a_valid & a_first_1;
	wire [1:0] _GEN_15 = (io_in_a_valid & a_first_1 ? 2'h1 : 2'h0);
	wire _T_1126 = a_first_done & a_first_1;
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? 4'h1 : 4'h0);
	wire [18:0] _a_opcodes_set_T_1 = {15'd0, a_opcodes_set_interm};
	wire [4:0] a_sizes_set_interm = (a_first_done & a_first_1 ? 5'h05 : 5'h00);
	wire [19:0] _a_sizes_set_T_1 = {15'd0, a_sizes_set_interm};
	wire _T_1130 = ~inflight;
	wire [1:0] _GEN_16 = (a_first_done & a_first_1 ? 2'h1 : 2'h0);
	wire [18:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [19:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 20'h00000);
	wire _T_1134 = io_in_d_valid & d_first_1;
	wire _T_1136 = ~_T_930;
	wire _T_1137 = (io_in_d_valid & d_first_1) & ~_T_930;
	wire [1:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_930 ? 2'h1 : 2'h0);
	wire [30:0] _d_opcodes_clr_T_5 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_sizes_clr_T_5 = {15'd0, _a_size_lookup_T_5};
	wire [30:0] _GEN_23 = (_T_1137 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [30:0] _GEN_24 = (_T_1137 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire _T_1149 = inflight | _T_1123;
	wire _T_1155 = _T_1007 | _T_1007;
	wire _T_1159 = 4'h2 == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1166 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1167 = (io_in_d_bits_opcode == _GEN_48) | _T_1166;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_75 = {4'd0, io_in_d_bits_size};
	wire _T_1171 = _GEN_75 == a_size_lookup;
	wire _T_1181 = ((_T_1134 & a_first_1) & io_in_a_valid) & _T_1136;
	wire a_set_wo_ready = _GEN_15[0];
	wire d_clr_wo_ready = _GEN_21[0];
	wire _T_1190 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire a_set = _GEN_16[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [7:0] a_sizes_set = _GEN_20[7:0];
	wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [7:0] d_sizes_clr = _GEN_24[7:0];
	wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1199 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [7:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [15:0] _GEN_78 = {8'd0, inflight_sizes_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_78 & _a_size_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_1225 = (io_in_d_valid & d_first_2) & _T_930;
	wire [30:0] _GEN_69 = (_T_1225 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1243 = _GEN_75 == c_size_lookup;
	wire [7:0] d_sizes_clr_1 = _GEN_69[7:0];
	wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 10'h000;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (io_in_d_valid)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (io_in_d_valid & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (io_in_d_valid & d_first)
			param_1 <= io_in_d_bits_param;
		if (io_in_d_valid & d_first)
			size_1 <= io_in_d_bits_size;
		if (io_in_d_valid & d_first)
			sink <= io_in_d_bits_sink;
		if (io_in_d_valid & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr_wo_ready;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 8'h00;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 10'h000;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (io_in_d_valid)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | io_in_d_valid)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 8'h00;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (io_in_d_valid)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module TLXbar_4 (
	clock,
	reset,
	auto_in_1_a_ready,
	auto_in_1_a_valid,
	auto_in_1_a_bits_address,
	auto_in_1_a_bits_data,
	auto_in_1_d_valid,
	auto_in_0_a_ready,
	auto_in_0_a_valid,
	auto_in_0_a_bits_opcode,
	auto_in_0_a_bits_param,
	auto_in_0_a_bits_size,
	auto_in_0_a_bits_source,
	auto_in_0_a_bits_address,
	auto_in_0_a_bits_mask,
	auto_in_0_a_bits_data,
	auto_in_0_a_bits_corrupt,
	auto_in_0_d_ready,
	auto_in_0_d_valid,
	auto_in_0_d_bits_opcode,
	auto_in_0_d_bits_param,
	auto_in_0_d_bits_size,
	auto_in_0_d_bits_source,
	auto_in_0_d_bits_sink,
	auto_in_0_d_bits_denied,
	auto_in_0_d_bits_data,
	auto_in_0_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_1_a_ready;
	input auto_in_1_a_valid;
	input [31:0] auto_in_1_a_bits_address;
	input [31:0] auto_in_1_a_bits_data;
	output wire auto_in_1_d_valid;
	output wire auto_in_0_a_ready;
	input auto_in_0_a_valid;
	input [2:0] auto_in_0_a_bits_opcode;
	input [2:0] auto_in_0_a_bits_param;
	input [3:0] auto_in_0_a_bits_size;
	input [1:0] auto_in_0_a_bits_source;
	input [31:0] auto_in_0_a_bits_address;
	input [3:0] auto_in_0_a_bits_mask;
	input [31:0] auto_in_0_a_bits_data;
	input auto_in_0_a_bits_corrupt;
	input auto_in_0_d_ready;
	output wire auto_in_0_d_valid;
	output wire [2:0] auto_in_0_d_bits_opcode;
	output wire [1:0] auto_in_0_d_bits_param;
	output wire [3:0] auto_in_0_d_bits_size;
	output wire [1:0] auto_in_0_d_bits_source;
	output wire auto_in_0_d_bits_sink;
	output wire auto_in_0_d_bits_denied;
	output wire [31:0] auto_in_0_d_bits_data;
	output wire auto_in_0_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire [1:0] monitor_io_in_a_bits_source;
	wire [31:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [3:0] monitor_io_in_d_bits_size;
	wire [1:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire monitor_1_clock;
	wire monitor_1_reset;
	wire monitor_1_io_in_a_ready;
	wire monitor_1_io_in_a_valid;
	wire [31:0] monitor_1_io_in_a_bits_address;
	wire monitor_1_io_in_d_valid;
	wire [2:0] monitor_1_io_in_d_bits_opcode;
	wire [1:0] monitor_1_io_in_d_bits_param;
	wire [3:0] monitor_1_io_in_d_bits_size;
	wire monitor_1_io_in_d_bits_sink;
	wire monitor_1_io_in_d_bits_denied;
	wire monitor_1_io_in_d_bits_corrupt;
	wire requestDOI_0_0 = ~auto_out_d_bits_source[2];
	wire requestDOI_0_1 = auto_out_d_bits_source == 3'h4;
	wire [26:0] _beatsAI_decode_T_1 = 27'h0000fff << auto_in_0_a_bits_size;
	wire [11:0] _beatsAI_decode_T_3 = ~_beatsAI_decode_T_1[11:0];
	wire [9:0] beatsAI_decode = _beatsAI_decode_T_3[11:2];
	wire beatsAI_opdata = ~auto_in_0_a_bits_opcode[2];
	reg [9:0] beatsLeft;
	wire idle = beatsLeft == 10'h000;
	wire latch = idle & auto_out_a_ready;
	wire [1:0] readys_valid = {auto_in_1_a_valid, auto_in_0_a_valid};
	wire _readys_T_3 = ~reset;
	reg [1:0] readys_mask;
	wire [1:0] _readys_filter_T = ~readys_mask;
	wire [1:0] _readys_filter_T_1 = readys_valid & _readys_filter_T;
	wire [3:0] readys_filter = {_readys_filter_T_1, auto_in_1_a_valid, auto_in_0_a_valid};
	wire [3:0] _GEN_1 = {1'd0, readys_filter[3:1]};
	wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_1;
	wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0};
	wire [3:0] _GEN_2 = {1'd0, _readys_unready_T_1[3:1]};
	wire [3:0] readys_unready = _GEN_2 | _readys_unready_T_4;
	wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0];
	wire [1:0] readys_readys = ~_readys_readys_T_2;
	wire [1:0] _readys_mask_T = readys_readys & readys_valid;
	wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0};
	wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0];
	wire readys_0 = readys_readys[0];
	wire readys_1 = readys_readys[1];
	wire earlyWinner_0 = readys_0 & auto_in_0_a_valid;
	wire earlyWinner_1 = readys_1 & auto_in_1_a_valid;
	wire _prefixOR_T = earlyWinner_0 | earlyWinner_1;
	wire _T_10 = auto_in_0_a_valid | auto_in_1_a_valid;
	wire _T_11 = ~(auto_in_0_a_valid | auto_in_1_a_valid);
	reg state_0;
	wire muxStateEarly_0 = (idle ? earlyWinner_0 : state_0);
	reg state_1;
	wire muxStateEarly_1 = (idle ? earlyWinner_1 : state_1);
	wire _out_0_a_earlyValid_T_3 = (state_0 & auto_in_0_a_valid) | (state_1 & auto_in_1_a_valid);
	wire out_2_0_a_earlyValid = (idle ? _T_10 : _out_0_a_earlyValid_T_3);
	wire _beatsLeft_T_2 = auto_out_a_ready & out_2_0_a_earlyValid;
	wire [9:0] _GEN_3 = {9'd0, _beatsLeft_T_2};
	wire [9:0] _beatsLeft_T_4 = beatsLeft - _GEN_3;
	wire allowed_0 = (idle ? readys_0 : state_0);
	wire allowed_1 = (idle ? readys_1 : state_1);
	wire [31:0] _T_27 = (muxStateEarly_0 ? auto_in_0_a_bits_data : 32'h00000000);
	wire [31:0] _T_28 = (muxStateEarly_1 ? auto_in_1_a_bits_data : 32'h00000000);
	wire [3:0] _T_30 = (muxStateEarly_0 ? auto_in_0_a_bits_mask : 4'h0);
	wire [3:0] _T_31 = (muxStateEarly_1 ? 4'hf : 4'h0);
	wire [31:0] _T_33 = (muxStateEarly_0 ? auto_in_0_a_bits_address : 32'h00000000);
	wire [31:0] _T_34 = (muxStateEarly_1 ? auto_in_1_a_bits_address : 32'h00000000);
	wire [2:0] in_0_a_bits_source = {1'd0, auto_in_0_a_bits_source};
	wire [2:0] _T_36 = (muxStateEarly_0 ? in_0_a_bits_source : 3'h0);
	wire [2:0] _T_37 = (muxStateEarly_1 ? 3'h4 : 3'h0);
	wire [3:0] _T_39 = (muxStateEarly_0 ? auto_in_0_a_bits_size : 4'h0);
	wire [3:0] _T_40 = (muxStateEarly_1 ? 4'h2 : 4'h0);
	TLMonitor_16 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	TLMonitor_17 monitor_1(
		.clock(monitor_1_clock),
		.reset(monitor_1_reset),
		.io_in_a_ready(monitor_1_io_in_a_ready),
		.io_in_a_valid(monitor_1_io_in_a_valid),
		.io_in_a_bits_address(monitor_1_io_in_a_bits_address),
		.io_in_d_valid(monitor_1_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_1_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_1_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_1_io_in_d_bits_size),
		.io_in_d_bits_sink(monitor_1_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_1_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_1_io_in_d_bits_corrupt)
	);
	assign auto_in_1_a_ready = auto_out_a_ready & allowed_1;
	assign auto_in_1_d_valid = auto_out_d_valid & requestDOI_0_1;
	assign auto_in_0_a_ready = auto_out_a_ready & allowed_0;
	assign auto_in_0_d_valid = auto_out_d_valid & requestDOI_0_0;
	assign auto_in_0_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_0_d_bits_param = auto_out_d_bits_param;
	assign auto_in_0_d_bits_size = auto_out_d_bits_size;
	assign auto_in_0_d_bits_source = auto_out_d_bits_source[1:0];
	assign auto_in_0_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_0_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_0_d_bits_data = auto_out_d_bits_data;
	assign auto_in_0_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = (idle ? _T_10 : _out_0_a_earlyValid_T_3);
	assign auto_out_a_bits_opcode = (muxStateEarly_0 ? auto_in_0_a_bits_opcode : 3'h0);
	assign auto_out_a_bits_param = (muxStateEarly_0 ? auto_in_0_a_bits_param : 3'h0);
	assign auto_out_a_bits_size = _T_39 | _T_40;
	assign auto_out_a_bits_source = _T_36 | _T_37;
	assign auto_out_a_bits_address = _T_33 | _T_34;
	assign auto_out_a_bits_mask = _T_30 | _T_31;
	assign auto_out_a_bits_data = _T_27 | _T_28;
	assign auto_out_a_bits_corrupt = muxStateEarly_0 & auto_in_0_a_bits_corrupt;
	assign auto_out_d_ready = (requestDOI_0_0 & auto_in_0_d_ready) | requestDOI_0_1;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_out_a_ready & allowed_0;
	assign monitor_io_in_a_valid = auto_in_0_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_0_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_0_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_0_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_0_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_0_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_0_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_0_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_0_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid & requestDOI_0_0;
	assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_io_in_d_bits_param = auto_out_d_bits_param;
	assign monitor_io_in_d_bits_size = auto_out_d_bits_size;
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source[1:0];
	assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink;
	assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied;
	assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign monitor_1_clock = clock;
	assign monitor_1_reset = reset;
	assign monitor_1_io_in_a_ready = auto_out_a_ready & allowed_1;
	assign monitor_1_io_in_a_valid = auto_in_1_a_valid;
	assign monitor_1_io_in_a_bits_address = auto_in_1_a_bits_address;
	assign monitor_1_io_in_d_valid = auto_out_d_valid & requestDOI_0_1;
	assign monitor_1_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_1_io_in_d_bits_param = auto_out_d_bits_param;
	assign monitor_1_io_in_d_bits_size = auto_out_d_bits_size;
	assign monitor_1_io_in_d_bits_sink = auto_out_d_bits_sink;
	assign monitor_1_io_in_d_bits_denied = auto_out_d_bits_denied;
	assign monitor_1_io_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	always @(posedge clock) begin
		if (reset)
			beatsLeft <= 10'h000;
		else if (latch) begin
			if (earlyWinner_0) begin
				if (beatsAI_opdata)
					beatsLeft <= beatsAI_decode;
				else
					beatsLeft <= 10'h000;
			end
			else
				beatsLeft <= 10'h000;
		end
		else
			beatsLeft <= _beatsLeft_T_4;
		if (reset)
			readys_mask <= 2'h3;
		else if (latch & |readys_valid)
			readys_mask <= _readys_mask_T_3;
		if (reset)
			state_0 <= 1'h0;
		else if (idle)
			state_0 <= earlyWinner_0;
		if (reset)
			state_1 <= 1'h0;
		else if (idle)
			state_1 <= earlyWinner_1;
	end
endmodule
module TLMonitor_18 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire _T_44 = io_in_a_bits_size <= 4'hc;
	wire _T_53 = _T_44 & source_ok;
	wire [32:0] _T_59 = $signed(_T_7) & -33'sh000005000;
	wire _T_60 = $signed(_T_59) == 33'sh000000000;
	wire [31:0] _T_61 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_62 = {1'b0, $signed(_T_61)};
	wire [32:0] _T_64 = $signed(_T_62) & -33'sh000001000;
	wire _T_65 = $signed(_T_64) == 33'sh000000000;
	wire [31:0] _T_66 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_67 = {1'b0, $signed(_T_66)};
	wire [32:0] _T_69 = $signed(_T_67) & -33'sh000010000;
	wire _T_70 = $signed(_T_69) == 33'sh000000000;
	wire [31:0] _T_71 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_72 = {1'b0, $signed(_T_71)};
	wire [32:0] _T_74 = $signed(_T_72) & -33'sh000010000;
	wire _T_75 = $signed(_T_74) == 33'sh000000000;
	wire [31:0] _T_76 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_77 = {1'b0, $signed(_T_76)};
	wire [32:0] _T_79 = $signed(_T_77) & -33'sh000011000;
	wire _T_80 = $signed(_T_79) == 33'sh000000000;
	wire [31:0] _T_81 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_82 = {1'b0, $signed(_T_81)};
	wire [32:0] _T_84 = $signed(_T_82) & -33'sh000010000;
	wire _T_85 = $signed(_T_84) == 33'sh000000000;
	wire [31:0] _T_86 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_87 = {1'b0, $signed(_T_86)};
	wire [32:0] _T_89 = $signed(_T_87) & -33'sh004000000;
	wire _T_90 = $signed(_T_89) == 33'sh000000000;
	wire [31:0] _T_91 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_92 = {1'b0, $signed(_T_91)};
	wire [32:0] _T_94 = $signed(_T_92) & -33'sh000001000;
	wire _T_95 = $signed(_T_94) == 33'sh000000000;
	wire [31:0] _T_96 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_97 = {1'b0, $signed(_T_96)};
	wire [32:0] _T_99 = $signed(_T_97) & -33'sh000001000;
	wire _T_100 = $signed(_T_99) == 33'sh000000000;
	wire [31:0] _T_101 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_102 = {1'b0, $signed(_T_101)};
	wire [32:0] _T_104 = $signed(_T_102) & -33'sh000004000;
	wire _T_105 = $signed(_T_104) == 33'sh000000000;
	wire _T_200 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_204 = ~io_in_a_bits_mask;
	wire _T_205 = _T_204 == 4'h0;
	wire _T_209 = ~io_in_a_bits_corrupt;
	wire _T_213 = io_in_a_bits_opcode == 3'h7;
	wire _T_375 = io_in_a_bits_param != 3'h0;
	wire _T_388 = io_in_a_bits_opcode == 3'h4;
	wire _T_413 = _T_44 & _T_65;
	wire _T_415 = io_in_a_bits_size <= 4'h6;
	wire _T_470 = (((((((_T_60 | _T_70) | _T_75) | _T_80) | _T_85) | _T_90) | _T_95) | _T_100) | _T_105;
	wire _T_471 = _T_415 & _T_470;
	wire _T_473 = _T_413 | _T_471;
	wire _T_483 = io_in_a_bits_param == 3'h0;
	wire _T_487 = io_in_a_bits_mask == mask;
	wire _T_495 = io_in_a_bits_opcode == 3'h0;
	wire _T_562 = (((((_T_60 | _T_80) | _T_85) | _T_90) | _T_95) | _T_100) | _T_105;
	wire _T_563 = _T_415 & _T_562;
	wire _T_578 = _T_413 | _T_563;
	wire _T_580 = _T_53 & _T_578;
	wire _T_598 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_697 = ~mask;
	wire [3:0] _T_698 = io_in_a_bits_mask & _T_697;
	wire _T_699 = _T_698 == 4'h0;
	wire _T_703 = io_in_a_bits_opcode == 3'h2;
	wire _T_717 = io_in_a_bits_size <= 4'h2;
	wire [31:0] _T_725 = io_in_a_bits_address ^ 32'h00004000;
	wire [32:0] _T_726 = {1'b0, $signed(_T_725)};
	wire [32:0] _T_728 = $signed(_T_726) & -33'sh000001000;
	wire _T_729 = $signed(_T_728) == 33'sh000000000;
	wire _T_742 = ((_T_65 | _T_729) | _T_95) | _T_100;
	wire _T_743 = _T_717 & _T_742;
	wire _T_781 = 4'h2 == io_in_a_bits_size;
	wire _T_788 = _T_781 & _T_105;
	wire _T_791 = _T_743 | _T_788;
	wire _T_792 = _T_53 & _T_791;
	wire _T_802 = io_in_a_bits_param <= 3'h4;
	wire _T_810 = io_in_a_bits_opcode == 3'h3;
	wire _T_909 = io_in_a_bits_param <= 3'h3;
	wire _T_917 = io_in_a_bits_opcode == 3'h5;
	wire _T_997 = _T_53 & _T_413;
	wire _T_1007 = io_in_a_bits_param <= 3'h1;
	wire _T_1019 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_1023 = io_in_d_bits_opcode == 3'h6;
	wire _T_1027 = io_in_d_bits_size >= 4'h2;
	wire _T_1031 = io_in_d_bits_param == 2'h0;
	wire _T_1035 = ~io_in_d_bits_corrupt;
	wire _T_1039 = ~io_in_d_bits_denied;
	wire _T_1043 = io_in_d_bits_opcode == 3'h4;
	wire _T_1054 = io_in_d_bits_param <= 2'h2;
	wire _T_1058 = io_in_d_bits_param != 2'h2;
	wire _T_1071 = io_in_d_bits_opcode == 3'h5;
	wire _T_1091 = _T_1039 | io_in_d_bits_corrupt;
	wire _T_1100 = io_in_d_bits_opcode == 3'h0;
	wire _T_1117 = io_in_d_bits_opcode == 3'h1;
	wire _T_1135 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg [2:0] source;
	reg [31:0] address;
	wire _T_1165 = io_in_a_valid & ~a_first;
	wire _T_1166 = io_in_a_bits_opcode == opcode;
	wire _T_1170 = io_in_a_bits_param == param;
	wire _T_1174 = io_in_a_bits_size == size;
	wire _T_1178 = io_in_a_bits_source == source;
	wire _T_1182 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_1189 = io_in_d_valid & ~d_first;
	wire _T_1190 = io_in_d_bits_opcode == opcode_1;
	wire _T_1194 = io_in_d_bits_param == param_1;
	wire _T_1198 = io_in_d_bits_size == size_1;
	wire _T_1202 = io_in_d_bits_source == source_1;
	wire _T_1206 = io_in_d_bits_sink == sink;
	wire _T_1210 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [39:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [5:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0};
	wire [39:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T;
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [39:0] _GEN_75 = {24'd0, _a_size_lookup_T_5};
	wire [39:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_75;
	wire [39:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[39:1]};
	wire _T_1216 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire _T_1219 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [4:0] _GEN_77 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_77};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [5:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [67:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [67:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire [4:0] _T_1221 = inflight >> io_in_a_bits_source;
	wire _T_1223 = ~_T_1221[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [67:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 68'h00000000000000000);
	wire _T_1227 = io_in_d_valid & d_first_1;
	wire _T_1229 = ~_T_1023;
	wire _T_1230 = (io_in_d_valid & d_first_1) & ~_T_1023;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [78:0] _GEN_4 = {63'd0, _a_size_lookup_T_5};
	wire [78:0] _d_sizes_clr_T_5 = _GEN_4 << _a_size_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_1229 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1229 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [78:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1229 ? _d_sizes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_1216 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_1240 = inflight >> io_in_d_bits_source;
	wire _T_1242 = _T_1240[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1247 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1248 = (io_in_d_bits_opcode == _GEN_32) | _T_1247;
	wire _T_1252 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1259 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1260 = (io_in_d_bits_opcode == _GEN_48) | _T_1259;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_79 = {4'd0, io_in_d_bits_size};
	wire _T_1264 = _GEN_79 == a_size_lookup;
	wire _T_1274 = (((_T_1227 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_1229;
	wire _T_1276 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [39:0] a_sizes_set = _GEN_20[39:0];
	wire [39:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [39:0] d_sizes_clr = _GEN_24[39:0];
	wire [39:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [39:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1285 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [39:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [39:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T;
	wire [39:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_75;
	wire [39:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[39:1]};
	wire _T_1311 = (io_in_d_valid & d_first_2) & _T_1023;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_1023 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_1023 ? _d_sizes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_1319 = inflight_1 >> io_in_d_bits_source;
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1329 = _GEN_79 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [39:0] d_sizes_clr_1 = _GEN_69[39:0];
	wire [39:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [39:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	reg [31:0] watchdog_1;
	wire _T_1349 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 40'h0000000000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 40'h0000000000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLXbar_5 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_8_a_ready,
	auto_out_8_a_valid,
	auto_out_8_a_bits_opcode,
	auto_out_8_a_bits_param,
	auto_out_8_a_bits_size,
	auto_out_8_a_bits_source,
	auto_out_8_a_bits_address,
	auto_out_8_a_bits_mask,
	auto_out_8_a_bits_data,
	auto_out_8_a_bits_corrupt,
	auto_out_8_d_ready,
	auto_out_8_d_valid,
	auto_out_8_d_bits_opcode,
	auto_out_8_d_bits_param,
	auto_out_8_d_bits_size,
	auto_out_8_d_bits_source,
	auto_out_8_d_bits_sink,
	auto_out_8_d_bits_denied,
	auto_out_8_d_bits_data,
	auto_out_8_d_bits_corrupt,
	auto_out_7_a_ready,
	auto_out_7_a_valid,
	auto_out_7_a_bits_opcode,
	auto_out_7_a_bits_param,
	auto_out_7_a_bits_size,
	auto_out_7_a_bits_source,
	auto_out_7_a_bits_address,
	auto_out_7_a_bits_mask,
	auto_out_7_a_bits_data,
	auto_out_7_a_bits_corrupt,
	auto_out_7_d_ready,
	auto_out_7_d_valid,
	auto_out_7_d_bits_opcode,
	auto_out_7_d_bits_param,
	auto_out_7_d_bits_size,
	auto_out_7_d_bits_source,
	auto_out_7_d_bits_sink,
	auto_out_7_d_bits_denied,
	auto_out_7_d_bits_data,
	auto_out_7_d_bits_corrupt,
	auto_out_6_a_ready,
	auto_out_6_a_valid,
	auto_out_6_a_bits_opcode,
	auto_out_6_a_bits_param,
	auto_out_6_a_bits_size,
	auto_out_6_a_bits_source,
	auto_out_6_a_bits_address,
	auto_out_6_a_bits_mask,
	auto_out_6_a_bits_corrupt,
	auto_out_6_d_ready,
	auto_out_6_d_valid,
	auto_out_6_d_bits_size,
	auto_out_6_d_bits_source,
	auto_out_6_d_bits_data,
	auto_out_5_a_ready,
	auto_out_5_a_valid,
	auto_out_5_a_bits_opcode,
	auto_out_5_a_bits_param,
	auto_out_5_a_bits_size,
	auto_out_5_a_bits_source,
	auto_out_5_a_bits_address,
	auto_out_5_a_bits_mask,
	auto_out_5_a_bits_data,
	auto_out_5_d_ready,
	auto_out_5_d_valid,
	auto_out_5_d_bits_opcode,
	auto_out_5_d_bits_param,
	auto_out_5_d_bits_size,
	auto_out_5_d_bits_source,
	auto_out_5_d_bits_sink,
	auto_out_5_d_bits_denied,
	auto_out_5_d_bits_data,
	auto_out_5_d_bits_corrupt,
	auto_out_4_a_ready,
	auto_out_4_a_valid,
	auto_out_4_a_bits_opcode,
	auto_out_4_a_bits_param,
	auto_out_4_a_bits_size,
	auto_out_4_a_bits_source,
	auto_out_4_a_bits_address,
	auto_out_4_a_bits_mask,
	auto_out_4_a_bits_data,
	auto_out_4_a_bits_corrupt,
	auto_out_4_d_ready,
	auto_out_4_d_valid,
	auto_out_4_d_bits_opcode,
	auto_out_4_d_bits_size,
	auto_out_4_d_bits_source,
	auto_out_4_d_bits_data,
	auto_out_3_a_ready,
	auto_out_3_a_valid,
	auto_out_3_a_bits_opcode,
	auto_out_3_a_bits_param,
	auto_out_3_a_bits_size,
	auto_out_3_a_bits_source,
	auto_out_3_a_bits_address,
	auto_out_3_a_bits_mask,
	auto_out_3_a_bits_data,
	auto_out_3_a_bits_corrupt,
	auto_out_3_d_ready,
	auto_out_3_d_valid,
	auto_out_3_d_bits_opcode,
	auto_out_3_d_bits_size,
	auto_out_3_d_bits_source,
	auto_out_3_d_bits_data,
	auto_out_2_a_ready,
	auto_out_2_a_valid,
	auto_out_2_a_bits_opcode,
	auto_out_2_a_bits_param,
	auto_out_2_a_bits_size,
	auto_out_2_a_bits_source,
	auto_out_2_a_bits_address,
	auto_out_2_a_bits_mask,
	auto_out_2_a_bits_data,
	auto_out_2_a_bits_corrupt,
	auto_out_2_d_ready,
	auto_out_2_d_valid,
	auto_out_2_d_bits_opcode,
	auto_out_2_d_bits_size,
	auto_out_2_d_bits_source,
	auto_out_2_d_bits_data,
	auto_out_1_a_ready,
	auto_out_1_a_valid,
	auto_out_1_a_bits_opcode,
	auto_out_1_a_bits_param,
	auto_out_1_a_bits_size,
	auto_out_1_a_bits_source,
	auto_out_1_a_bits_address,
	auto_out_1_a_bits_mask,
	auto_out_1_a_bits_data,
	auto_out_1_a_bits_corrupt,
	auto_out_1_d_ready,
	auto_out_1_d_valid,
	auto_out_1_d_bits_opcode,
	auto_out_1_d_bits_param,
	auto_out_1_d_bits_size,
	auto_out_1_d_bits_source,
	auto_out_1_d_bits_sink,
	auto_out_1_d_bits_denied,
	auto_out_1_d_bits_data,
	auto_out_1_d_bits_corrupt,
	auto_out_0_a_ready,
	auto_out_0_a_valid,
	auto_out_0_a_bits_opcode,
	auto_out_0_a_bits_param,
	auto_out_0_a_bits_size,
	auto_out_0_a_bits_source,
	auto_out_0_a_bits_address,
	auto_out_0_a_bits_mask,
	auto_out_0_a_bits_corrupt,
	auto_out_0_d_ready,
	auto_out_0_d_valid,
	auto_out_0_d_bits_opcode,
	auto_out_0_d_bits_param,
	auto_out_0_d_bits_size,
	auto_out_0_d_bits_source,
	auto_out_0_d_bits_sink,
	auto_out_0_d_bits_denied,
	auto_out_0_d_bits_data,
	auto_out_0_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_8_a_ready;
	output wire auto_out_8_a_valid;
	output wire [2:0] auto_out_8_a_bits_opcode;
	output wire [2:0] auto_out_8_a_bits_param;
	output wire [2:0] auto_out_8_a_bits_size;
	output wire [2:0] auto_out_8_a_bits_source;
	output wire [20:0] auto_out_8_a_bits_address;
	output wire [3:0] auto_out_8_a_bits_mask;
	output wire [31:0] auto_out_8_a_bits_data;
	output wire auto_out_8_a_bits_corrupt;
	output wire auto_out_8_d_ready;
	input auto_out_8_d_valid;
	input [2:0] auto_out_8_d_bits_opcode;
	input [1:0] auto_out_8_d_bits_param;
	input [2:0] auto_out_8_d_bits_size;
	input [2:0] auto_out_8_d_bits_source;
	input auto_out_8_d_bits_sink;
	input auto_out_8_d_bits_denied;
	input [31:0] auto_out_8_d_bits_data;
	input auto_out_8_d_bits_corrupt;
	input auto_out_7_a_ready;
	output wire auto_out_7_a_valid;
	output wire [2:0] auto_out_7_a_bits_opcode;
	output wire [2:0] auto_out_7_a_bits_param;
	output wire [2:0] auto_out_7_a_bits_size;
	output wire [2:0] auto_out_7_a_bits_source;
	output wire [20:0] auto_out_7_a_bits_address;
	output wire [3:0] auto_out_7_a_bits_mask;
	output wire [31:0] auto_out_7_a_bits_data;
	output wire auto_out_7_a_bits_corrupt;
	output wire auto_out_7_d_ready;
	input auto_out_7_d_valid;
	input [2:0] auto_out_7_d_bits_opcode;
	input [1:0] auto_out_7_d_bits_param;
	input [2:0] auto_out_7_d_bits_size;
	input [2:0] auto_out_7_d_bits_source;
	input auto_out_7_d_bits_sink;
	input auto_out_7_d_bits_denied;
	input [31:0] auto_out_7_d_bits_data;
	input auto_out_7_d_bits_corrupt;
	input auto_out_6_a_ready;
	output wire auto_out_6_a_valid;
	output wire [2:0] auto_out_6_a_bits_opcode;
	output wire [2:0] auto_out_6_a_bits_param;
	output wire [2:0] auto_out_6_a_bits_size;
	output wire [2:0] auto_out_6_a_bits_source;
	output wire [16:0] auto_out_6_a_bits_address;
	output wire [3:0] auto_out_6_a_bits_mask;
	output wire auto_out_6_a_bits_corrupt;
	output wire auto_out_6_d_ready;
	input auto_out_6_d_valid;
	input [2:0] auto_out_6_d_bits_size;
	input [2:0] auto_out_6_d_bits_source;
	input [31:0] auto_out_6_d_bits_data;
	input auto_out_5_a_ready;
	output wire auto_out_5_a_valid;
	output wire [2:0] auto_out_5_a_bits_opcode;
	output wire [2:0] auto_out_5_a_bits_param;
	output wire [2:0] auto_out_5_a_bits_size;
	output wire [2:0] auto_out_5_a_bits_source;
	output wire [31:0] auto_out_5_a_bits_address;
	output wire [3:0] auto_out_5_a_bits_mask;
	output wire [31:0] auto_out_5_a_bits_data;
	output wire auto_out_5_d_ready;
	input auto_out_5_d_valid;
	input [2:0] auto_out_5_d_bits_opcode;
	input [1:0] auto_out_5_d_bits_param;
	input [2:0] auto_out_5_d_bits_size;
	input [2:0] auto_out_5_d_bits_source;
	input auto_out_5_d_bits_sink;
	input auto_out_5_d_bits_denied;
	input [31:0] auto_out_5_d_bits_data;
	input auto_out_5_d_bits_corrupt;
	input auto_out_4_a_ready;
	output wire auto_out_4_a_valid;
	output wire [2:0] auto_out_4_a_bits_opcode;
	output wire [2:0] auto_out_4_a_bits_param;
	output wire [2:0] auto_out_4_a_bits_size;
	output wire [2:0] auto_out_4_a_bits_source;
	output wire [11:0] auto_out_4_a_bits_address;
	output wire [3:0] auto_out_4_a_bits_mask;
	output wire [31:0] auto_out_4_a_bits_data;
	output wire auto_out_4_a_bits_corrupt;
	output wire auto_out_4_d_ready;
	input auto_out_4_d_valid;
	input [2:0] auto_out_4_d_bits_opcode;
	input [2:0] auto_out_4_d_bits_size;
	input [2:0] auto_out_4_d_bits_source;
	input [31:0] auto_out_4_d_bits_data;
	input auto_out_3_a_ready;
	output wire auto_out_3_a_valid;
	output wire [2:0] auto_out_3_a_bits_opcode;
	output wire [2:0] auto_out_3_a_bits_param;
	output wire [2:0] auto_out_3_a_bits_size;
	output wire [2:0] auto_out_3_a_bits_source;
	output wire [25:0] auto_out_3_a_bits_address;
	output wire [3:0] auto_out_3_a_bits_mask;
	output wire [31:0] auto_out_3_a_bits_data;
	output wire auto_out_3_a_bits_corrupt;
	output wire auto_out_3_d_ready;
	input auto_out_3_d_valid;
	input [2:0] auto_out_3_d_bits_opcode;
	input [2:0] auto_out_3_d_bits_size;
	input [2:0] auto_out_3_d_bits_source;
	input [31:0] auto_out_3_d_bits_data;
	input auto_out_2_a_ready;
	output wire auto_out_2_a_valid;
	output wire [2:0] auto_out_2_a_bits_opcode;
	output wire [2:0] auto_out_2_a_bits_param;
	output wire [2:0] auto_out_2_a_bits_size;
	output wire [2:0] auto_out_2_a_bits_source;
	output wire [27:0] auto_out_2_a_bits_address;
	output wire [3:0] auto_out_2_a_bits_mask;
	output wire [31:0] auto_out_2_a_bits_data;
	output wire auto_out_2_a_bits_corrupt;
	output wire auto_out_2_d_ready;
	input auto_out_2_d_valid;
	input [2:0] auto_out_2_d_bits_opcode;
	input [2:0] auto_out_2_d_bits_size;
	input [2:0] auto_out_2_d_bits_source;
	input [31:0] auto_out_2_d_bits_data;
	input auto_out_1_a_ready;
	output wire auto_out_1_a_valid;
	output wire [2:0] auto_out_1_a_bits_opcode;
	output wire [2:0] auto_out_1_a_bits_param;
	output wire [2:0] auto_out_1_a_bits_size;
	output wire [2:0] auto_out_1_a_bits_source;
	output wire [30:0] auto_out_1_a_bits_address;
	output wire [3:0] auto_out_1_a_bits_mask;
	output wire [31:0] auto_out_1_a_bits_data;
	output wire auto_out_1_a_bits_corrupt;
	output wire auto_out_1_d_ready;
	input auto_out_1_d_valid;
	input [2:0] auto_out_1_d_bits_opcode;
	input [1:0] auto_out_1_d_bits_param;
	input [2:0] auto_out_1_d_bits_size;
	input [2:0] auto_out_1_d_bits_source;
	input auto_out_1_d_bits_sink;
	input auto_out_1_d_bits_denied;
	input [31:0] auto_out_1_d_bits_data;
	input auto_out_1_d_bits_corrupt;
	input auto_out_0_a_ready;
	output wire auto_out_0_a_valid;
	output wire [2:0] auto_out_0_a_bits_opcode;
	output wire [2:0] auto_out_0_a_bits_param;
	output wire [3:0] auto_out_0_a_bits_size;
	output wire [2:0] auto_out_0_a_bits_source;
	output wire [13:0] auto_out_0_a_bits_address;
	output wire [3:0] auto_out_0_a_bits_mask;
	output wire auto_out_0_a_bits_corrupt;
	output wire auto_out_0_d_ready;
	input auto_out_0_d_valid;
	input [2:0] auto_out_0_d_bits_opcode;
	input [1:0] auto_out_0_d_bits_param;
	input [3:0] auto_out_0_d_bits_size;
	input [2:0] auto_out_0_d_bits_source;
	input auto_out_0_d_bits_sink;
	input auto_out_0_d_bits_denied;
	input [31:0] auto_out_0_d_bits_data;
	input auto_out_0_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [31:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [3:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	reg [9:0] beatsLeft;
	wire idle = beatsLeft == 10'h000;
	wire [8:0] readys_valid = {auto_out_8_d_valid, auto_out_7_d_valid, auto_out_6_d_valid, auto_out_5_d_valid, auto_out_4_d_valid, auto_out_3_d_valid, auto_out_2_d_valid, auto_out_1_d_valid, auto_out_0_d_valid};
	reg [8:0] readys_mask;
	wire [8:0] _readys_filter_T = ~readys_mask;
	wire [8:0] _readys_filter_T_1 = readys_valid & _readys_filter_T;
	wire [17:0] readys_filter = {_readys_filter_T_1, auto_out_8_d_valid, auto_out_7_d_valid, auto_out_6_d_valid, auto_out_5_d_valid, auto_out_4_d_valid, auto_out_3_d_valid, auto_out_2_d_valid, auto_out_1_d_valid, auto_out_0_d_valid};
	wire [17:0] _GEN_1 = {1'd0, readys_filter[17:1]};
	wire [17:0] _readys_unready_T_1 = readys_filter | _GEN_1;
	wire [17:0] _GEN_2 = {2'd0, _readys_unready_T_1[17:2]};
	wire [17:0] _readys_unready_T_3 = _readys_unready_T_1 | _GEN_2;
	wire [17:0] _GEN_3 = {4'd0, _readys_unready_T_3[17:4]};
	wire [17:0] _readys_unready_T_5 = _readys_unready_T_3 | _GEN_3;
	wire [17:0] _GEN_4 = {8'd0, _readys_unready_T_5[17:8]};
	wire [17:0] _readys_unready_T_7 = _readys_unready_T_5 | _GEN_4;
	wire [17:0] _readys_unready_T_10 = {readys_mask, 9'h000};
	wire [17:0] _GEN_5 = {1'd0, _readys_unready_T_7[17:1]};
	wire [17:0] readys_unready = _GEN_5 | _readys_unready_T_10;
	wire [8:0] _readys_readys_T_2 = readys_unready[17:9] & readys_unready[8:0];
	wire [8:0] readys_readys = ~_readys_readys_T_2;
	wire readys_0 = readys_readys[0];
	wire earlyWinner_0 = readys_0 & auto_out_0_d_valid;
	reg state_0;
	wire muxStateEarly_0 = (idle ? earlyWinner_0 : state_0);
	wire [2:0] _T_148 = (muxStateEarly_0 ? auto_out_0_d_bits_source : 3'h0);
	wire readys_1 = readys_readys[1];
	wire earlyWinner_1 = readys_1 & auto_out_1_d_valid;
	reg state_1;
	wire muxStateEarly_1 = (idle ? earlyWinner_1 : state_1);
	wire [2:0] _T_149 = (muxStateEarly_1 ? auto_out_1_d_bits_source : 3'h0);
	wire [2:0] _T_157 = _T_148 | _T_149;
	wire readys_2 = readys_readys[2];
	wire earlyWinner_2 = readys_2 & auto_out_2_d_valid;
	reg state_2;
	wire muxStateEarly_2 = (idle ? earlyWinner_2 : state_2);
	wire [2:0] _T_150 = (muxStateEarly_2 ? auto_out_2_d_bits_source : 3'h0);
	wire [2:0] _T_158 = _T_157 | _T_150;
	wire readys_3 = readys_readys[3];
	wire earlyWinner_3 = readys_3 & auto_out_3_d_valid;
	reg state_3;
	wire muxStateEarly_3 = (idle ? earlyWinner_3 : state_3);
	wire [2:0] _T_151 = (muxStateEarly_3 ? auto_out_3_d_bits_source : 3'h0);
	wire [2:0] _T_159 = _T_158 | _T_151;
	wire readys_4 = readys_readys[4];
	wire earlyWinner_4 = readys_4 & auto_out_4_d_valid;
	reg state_4;
	wire muxStateEarly_4 = (idle ? earlyWinner_4 : state_4);
	wire [2:0] _T_152 = (muxStateEarly_4 ? auto_out_4_d_bits_source : 3'h0);
	wire [2:0] _T_160 = _T_159 | _T_152;
	wire readys_5 = readys_readys[5];
	wire earlyWinner_5 = readys_5 & auto_out_5_d_valid;
	reg state_5;
	wire muxStateEarly_5 = (idle ? earlyWinner_5 : state_5);
	wire [2:0] _T_153 = (muxStateEarly_5 ? auto_out_5_d_bits_source : 3'h0);
	wire [2:0] _T_161 = _T_160 | _T_153;
	wire readys_6 = readys_readys[6];
	wire earlyWinner_6 = readys_6 & auto_out_6_d_valid;
	reg state_6;
	wire muxStateEarly_6 = (idle ? earlyWinner_6 : state_6);
	wire [2:0] _T_154 = (muxStateEarly_6 ? auto_out_6_d_bits_source : 3'h0);
	wire [2:0] _T_162 = _T_161 | _T_154;
	wire readys_7 = readys_readys[7];
	wire earlyWinner_7 = readys_7 & auto_out_7_d_valid;
	reg state_7;
	wire muxStateEarly_7 = (idle ? earlyWinner_7 : state_7);
	wire [2:0] _T_155 = (muxStateEarly_7 ? auto_out_7_d_bits_source : 3'h0);
	wire [2:0] _T_163 = _T_162 | _T_155;
	wire readys_8 = readys_readys[8];
	wire earlyWinner_8 = readys_8 & auto_out_8_d_valid;
	reg state_8;
	wire muxStateEarly_8 = (idle ? earlyWinner_8 : state_8);
	wire [2:0] _T_156 = (muxStateEarly_8 ? auto_out_8_d_bits_source : 3'h0);
	wire [31:0] _requestAIO_T = auto_in_a_bits_address ^ 32'h00002000;
	wire [32:0] _requestAIO_T_1 = {1'b0, $signed(_requestAIO_T)};
	wire [32:0] _requestAIO_T_3 = $signed(_requestAIO_T_1) & 33'sh096136000;
	wire requestAIO_0_0 = $signed(_requestAIO_T_3) == 33'sh000000000;
	wire [31:0] _requestAIO_T_5 = auto_in_a_bits_address ^ 32'h00004000;
	wire [32:0] _requestAIO_T_6 = {1'b0, $signed(_requestAIO_T_5)};
	wire [32:0] _requestAIO_T_8 = $signed(_requestAIO_T_6) & 33'sh096136000;
	wire _requestAIO_T_9 = $signed(_requestAIO_T_8) == 33'sh000000000;
	wire [31:0] _requestAIO_T_10 = auto_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _requestAIO_T_11 = {1'b0, $signed(_requestAIO_T_10)};
	wire [32:0] _requestAIO_T_13 = $signed(_requestAIO_T_11) & 33'sh096130000;
	wire _requestAIO_T_14 = $signed(_requestAIO_T_13) == 33'sh000000000;
	wire [31:0] _requestAIO_T_15 = auto_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _requestAIO_T_16 = {1'b0, $signed(_requestAIO_T_15)};
	wire [32:0] _requestAIO_T_18 = $signed(_requestAIO_T_16) & 33'sh092136000;
	wire _requestAIO_T_19 = $signed(_requestAIO_T_18) == 33'sh000000000;
	wire requestAIO_0_1 = (_requestAIO_T_9 | _requestAIO_T_14) | _requestAIO_T_19;
	wire [31:0] _requestAIO_T_22 = auto_in_a_bits_address ^ 32'h04000000;
	wire [32:0] _requestAIO_T_23 = {1'b0, $signed(_requestAIO_T_22)};
	wire [32:0] _requestAIO_T_25 = $signed(_requestAIO_T_23) & 33'sh094000000;
	wire requestAIO_0_2 = $signed(_requestAIO_T_25) == 33'sh000000000;
	wire [31:0] _requestAIO_T_27 = auto_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _requestAIO_T_28 = {1'b0, $signed(_requestAIO_T_27)};
	wire [32:0] _requestAIO_T_30 = $signed(_requestAIO_T_28) & 33'sh096130000;
	wire requestAIO_0_3 = $signed(_requestAIO_T_30) == 33'sh000000000;
	wire [32:0] _requestAIO_T_33 = {1'b0, $signed(auto_in_a_bits_address)};
	wire [32:0] _requestAIO_T_35 = $signed(_requestAIO_T_33) & 33'sh096136000;
	wire requestAIO_0_4 = $signed(_requestAIO_T_35) == 33'sh000000000;
	wire [31:0] _requestAIO_T_37 = auto_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _requestAIO_T_38 = {1'b0, $signed(_requestAIO_T_37)};
	wire [32:0] _requestAIO_T_40 = $signed(_requestAIO_T_38) & 33'sh096134000;
	wire requestAIO_0_5 = $signed(_requestAIO_T_40) == 33'sh000000000;
	wire [31:0] _requestAIO_T_42 = auto_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _requestAIO_T_43 = {1'b0, $signed(_requestAIO_T_42)};
	wire [32:0] _requestAIO_T_45 = $signed(_requestAIO_T_43) & 33'sh096130000;
	wire requestAIO_0_6 = $signed(_requestAIO_T_45) == 33'sh000000000;
	wire [31:0] _requestAIO_T_47 = auto_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _requestAIO_T_48 = {1'b0, $signed(_requestAIO_T_47)};
	wire [32:0] _requestAIO_T_50 = $signed(_requestAIO_T_48) & 33'sh096136000;
	wire requestAIO_0_7 = $signed(_requestAIO_T_50) == 33'sh000000000;
	wire [31:0] _requestAIO_T_52 = auto_in_a_bits_address ^ 32'h00110000;
	wire [32:0] _requestAIO_T_53 = {1'b0, $signed(_requestAIO_T_52)};
	wire [32:0] _requestAIO_T_55 = $signed(_requestAIO_T_53) & 33'sh096136000;
	wire requestAIO_0_8 = $signed(_requestAIO_T_55) == 33'sh000000000;
	wire [26:0] _beatsDO_decode_T_1 = 27'h0000fff << auto_out_0_d_bits_size;
	wire [11:0] _beatsDO_decode_T_3 = ~_beatsDO_decode_T_1[11:0];
	wire [9:0] beatsDO_decode = _beatsDO_decode_T_3[11:2];
	wire beatsDO_opdata = auto_out_0_d_bits_opcode[0];
	wire [9:0] beatsDO_0 = (beatsDO_opdata ? beatsDO_decode : 10'h000);
	wire [3:0] out_1_1_d_bits_size = {1'd0, auto_out_1_d_bits_size};
	wire [20:0] _beatsDO_decode_T_5 = 21'h00003f << out_1_1_d_bits_size;
	wire [5:0] _beatsDO_decode_T_7 = ~_beatsDO_decode_T_5[5:0];
	wire [3:0] beatsDO_decode_1 = _beatsDO_decode_T_7[5:2];
	wire beatsDO_opdata_1 = auto_out_1_d_bits_opcode[0];
	wire [3:0] beatsDO_1 = (beatsDO_opdata_1 ? beatsDO_decode_1 : 4'h0);
	wire [3:0] out_1_2_d_bits_size = {1'd0, auto_out_2_d_bits_size};
	wire [20:0] _beatsDO_decode_T_9 = 21'h00003f << out_1_2_d_bits_size;
	wire [5:0] _beatsDO_decode_T_11 = ~_beatsDO_decode_T_9[5:0];
	wire [3:0] beatsDO_decode_2 = _beatsDO_decode_T_11[5:2];
	wire beatsDO_opdata_2 = auto_out_2_d_bits_opcode[0];
	wire [3:0] beatsDO_2 = (beatsDO_opdata_2 ? beatsDO_decode_2 : 4'h0);
	wire [3:0] out_1_3_d_bits_size = {1'd0, auto_out_3_d_bits_size};
	wire [20:0] _beatsDO_decode_T_13 = 21'h00003f << out_1_3_d_bits_size;
	wire [5:0] _beatsDO_decode_T_15 = ~_beatsDO_decode_T_13[5:0];
	wire [3:0] beatsDO_decode_3 = _beatsDO_decode_T_15[5:2];
	wire beatsDO_opdata_3 = auto_out_3_d_bits_opcode[0];
	wire [3:0] beatsDO_3 = (beatsDO_opdata_3 ? beatsDO_decode_3 : 4'h0);
	wire [3:0] out_1_4_d_bits_size = {1'd0, auto_out_4_d_bits_size};
	wire [20:0] _beatsDO_decode_T_17 = 21'h00003f << out_1_4_d_bits_size;
	wire [5:0] _beatsDO_decode_T_19 = ~_beatsDO_decode_T_17[5:0];
	wire [3:0] beatsDO_decode_4 = _beatsDO_decode_T_19[5:2];
	wire beatsDO_opdata_4 = auto_out_4_d_bits_opcode[0];
	wire [3:0] beatsDO_4 = (beatsDO_opdata_4 ? beatsDO_decode_4 : 4'h0);
	wire [3:0] out_1_5_d_bits_size = {1'd0, auto_out_5_d_bits_size};
	wire [20:0] _beatsDO_decode_T_21 = 21'h00003f << out_1_5_d_bits_size;
	wire [5:0] _beatsDO_decode_T_23 = ~_beatsDO_decode_T_21[5:0];
	wire [3:0] beatsDO_decode_5 = _beatsDO_decode_T_23[5:2];
	wire beatsDO_opdata_5 = auto_out_5_d_bits_opcode[0];
	wire [3:0] beatsDO_5 = (beatsDO_opdata_5 ? beatsDO_decode_5 : 4'h0);
	wire [3:0] out_1_6_d_bits_size = {1'd0, auto_out_6_d_bits_size};
	wire [20:0] _beatsDO_decode_T_25 = 21'h00003f << out_1_6_d_bits_size;
	wire [5:0] _beatsDO_decode_T_27 = ~_beatsDO_decode_T_25[5:0];
	wire [3:0] beatsDO_decode_6 = _beatsDO_decode_T_27[5:2];
	wire [3:0] out_1_7_d_bits_size = {1'd0, auto_out_7_d_bits_size};
	wire [20:0] _beatsDO_decode_T_29 = 21'h00003f << out_1_7_d_bits_size;
	wire [5:0] _beatsDO_decode_T_31 = ~_beatsDO_decode_T_29[5:0];
	wire [3:0] beatsDO_decode_7 = _beatsDO_decode_T_31[5:2];
	wire beatsDO_opdata_7 = auto_out_7_d_bits_opcode[0];
	wire [3:0] beatsDO_7 = (beatsDO_opdata_7 ? beatsDO_decode_7 : 4'h0);
	wire [3:0] out_1_8_d_bits_size = {1'd0, auto_out_8_d_bits_size};
	wire [20:0] _beatsDO_decode_T_33 = 21'h00003f << out_1_8_d_bits_size;
	wire [5:0] _beatsDO_decode_T_35 = ~_beatsDO_decode_T_33[5:0];
	wire [3:0] beatsDO_decode_8 = _beatsDO_decode_T_35[5:2];
	wire beatsDO_opdata_8 = auto_out_8_d_bits_opcode[0];
	wire [3:0] beatsDO_8 = (beatsDO_opdata_8 ? beatsDO_decode_8 : 4'h0);
	wire latch = idle & auto_in_d_ready;
	wire _readys_T_3 = ~reset;
	wire [8:0] _readys_mask_T = readys_readys & readys_valid;
	wire [9:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0};
	wire [8:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[8:0];
	wire [10:0] _readys_mask_T_4 = {_readys_mask_T_3, 2'h0};
	wire [8:0] _readys_mask_T_6 = _readys_mask_T_3 | _readys_mask_T_4[8:0];
	wire [12:0] _readys_mask_T_7 = {_readys_mask_T_6, 4'h0};
	wire [8:0] _readys_mask_T_9 = _readys_mask_T_6 | _readys_mask_T_7[8:0];
	wire [16:0] _readys_mask_T_10 = {_readys_mask_T_9, 8'h00};
	wire [8:0] _readys_mask_T_12 = _readys_mask_T_9 | _readys_mask_T_10[8:0];
	wire prefixOR_2 = earlyWinner_0 | earlyWinner_1;
	wire prefixOR_3 = prefixOR_2 | earlyWinner_2;
	wire prefixOR_4 = prefixOR_3 | earlyWinner_3;
	wire prefixOR_5 = prefixOR_4 | earlyWinner_4;
	wire prefixOR_6 = prefixOR_5 | earlyWinner_5;
	wire prefixOR_7 = prefixOR_6 | earlyWinner_6;
	wire prefixOR_8 = prefixOR_7 | earlyWinner_7;
	wire _prefixOR_T = prefixOR_8 | earlyWinner_8;
	wire _T_26 = ~prefixOR_8 | ~earlyWinner_8;
	wire _T_45 = (((((((auto_out_0_d_valid | auto_out_1_d_valid) | auto_out_2_d_valid) | auto_out_3_d_valid) | auto_out_4_d_valid) | auto_out_5_d_valid) | auto_out_6_d_valid) | auto_out_7_d_valid) | auto_out_8_d_valid;
	wire _T_46 = ~((((((((auto_out_0_d_valid | auto_out_1_d_valid) | auto_out_2_d_valid) | auto_out_3_d_valid) | auto_out_4_d_valid) | auto_out_5_d_valid) | auto_out_6_d_valid) | auto_out_7_d_valid) | auto_out_8_d_valid);
	wire [9:0] maskedBeats_0 = (earlyWinner_0 ? beatsDO_0 : 10'h000);
	wire [3:0] maskedBeats_1 = (earlyWinner_1 ? beatsDO_1 : 4'h0);
	wire [3:0] maskedBeats_2 = (earlyWinner_2 ? beatsDO_2 : 4'h0);
	wire [3:0] maskedBeats_3 = (earlyWinner_3 ? beatsDO_3 : 4'h0);
	wire [3:0] maskedBeats_4 = (earlyWinner_4 ? beatsDO_4 : 4'h0);
	wire [3:0] maskedBeats_5 = (earlyWinner_5 ? beatsDO_5 : 4'h0);
	wire [3:0] maskedBeats_6 = (earlyWinner_6 ? beatsDO_decode_6 : 4'h0);
	wire [3:0] maskedBeats_7 = (earlyWinner_7 ? beatsDO_7 : 4'h0);
	wire [3:0] maskedBeats_8 = (earlyWinner_8 ? beatsDO_8 : 4'h0);
	wire [9:0] _GEN_6 = {6'd0, maskedBeats_1};
	wire [9:0] _initBeats_T = maskedBeats_0 | _GEN_6;
	wire [9:0] _GEN_7 = {6'd0, maskedBeats_2};
	wire [9:0] _initBeats_T_1 = _initBeats_T | _GEN_7;
	wire [9:0] _GEN_8 = {6'd0, maskedBeats_3};
	wire [9:0] _initBeats_T_2 = _initBeats_T_1 | _GEN_8;
	wire [9:0] _GEN_9 = {6'd0, maskedBeats_4};
	wire [9:0] _initBeats_T_3 = _initBeats_T_2 | _GEN_9;
	wire [9:0] _GEN_10 = {6'd0, maskedBeats_5};
	wire [9:0] _initBeats_T_4 = _initBeats_T_3 | _GEN_10;
	wire [9:0] _GEN_11 = {6'd0, maskedBeats_6};
	wire [9:0] _initBeats_T_5 = _initBeats_T_4 | _GEN_11;
	wire [9:0] _GEN_12 = {6'd0, maskedBeats_7};
	wire [9:0] _initBeats_T_6 = _initBeats_T_5 | _GEN_12;
	wire [9:0] _GEN_13 = {6'd0, maskedBeats_8};
	wire [9:0] initBeats = _initBeats_T_6 | _GEN_13;
	wire _sink_ACancel_earlyValid_T_24 = ((((((((state_0 & auto_out_0_d_valid) | (state_1 & auto_out_1_d_valid)) | (state_2 & auto_out_2_d_valid)) | (state_3 & auto_out_3_d_valid)) | (state_4 & auto_out_4_d_valid)) | (state_5 & auto_out_5_d_valid)) | (state_6 & auto_out_6_d_valid)) | (state_7 & auto_out_7_d_valid)) | (state_8 & auto_out_8_d_valid);
	wire sink_ACancel_19_earlyValid = (idle ? _T_45 : _sink_ACancel_earlyValid_T_24);
	wire _beatsLeft_T_2 = auto_in_d_ready & sink_ACancel_19_earlyValid;
	wire [9:0] _GEN_14 = {9'd0, _beatsLeft_T_2};
	wire [9:0] _beatsLeft_T_4 = beatsLeft - _GEN_14;
	wire allowed_0 = (idle ? readys_0 : state_0);
	wire allowed_1 = (idle ? readys_1 : state_1);
	wire allowed_2 = (idle ? readys_2 : state_2);
	wire allowed_3 = (idle ? readys_3 : state_3);
	wire allowed_4 = (idle ? readys_4 : state_4);
	wire allowed_5 = (idle ? readys_5 : state_5);
	wire allowed_6 = (idle ? readys_6 : state_6);
	wire allowed_7 = (idle ? readys_7 : state_7);
	wire allowed_8 = (idle ? readys_8 : state_8);
	wire [31:0] _T_97 = (muxStateEarly_0 ? auto_out_0_d_bits_data : 32'h00000000);
	wire [31:0] _T_98 = (muxStateEarly_1 ? auto_out_1_d_bits_data : 32'h00000000);
	wire [31:0] _T_99 = (muxStateEarly_2 ? auto_out_2_d_bits_data : 32'h00000000);
	wire [31:0] _T_100 = (muxStateEarly_3 ? auto_out_3_d_bits_data : 32'h00000000);
	wire [31:0] _T_101 = (muxStateEarly_4 ? auto_out_4_d_bits_data : 32'h00000000);
	wire [31:0] _T_102 = (muxStateEarly_5 ? auto_out_5_d_bits_data : 32'h00000000);
	wire [31:0] _T_103 = (muxStateEarly_6 ? auto_out_6_d_bits_data : 32'h00000000);
	wire [31:0] _T_104 = (muxStateEarly_7 ? auto_out_7_d_bits_data : 32'h00000000);
	wire [31:0] _T_105 = (muxStateEarly_8 ? auto_out_8_d_bits_data : 32'h00000000);
	wire [31:0] _T_106 = _T_97 | _T_98;
	wire [31:0] _T_107 = _T_106 | _T_99;
	wire [31:0] _T_108 = _T_107 | _T_100;
	wire [31:0] _T_109 = _T_108 | _T_101;
	wire [31:0] _T_110 = _T_109 | _T_102;
	wire [31:0] _T_111 = _T_110 | _T_103;
	wire [31:0] _T_112 = _T_111 | _T_104;
	wire [3:0] _T_165 = (muxStateEarly_0 ? auto_out_0_d_bits_size : 4'h0);
	wire [3:0] _T_166 = (muxStateEarly_1 ? out_1_1_d_bits_size : 4'h0);
	wire [3:0] _T_167 = (muxStateEarly_2 ? out_1_2_d_bits_size : 4'h0);
	wire [3:0] _T_168 = (muxStateEarly_3 ? out_1_3_d_bits_size : 4'h0);
	wire [3:0] _T_169 = (muxStateEarly_4 ? out_1_4_d_bits_size : 4'h0);
	wire [3:0] _T_170 = (muxStateEarly_5 ? out_1_5_d_bits_size : 4'h0);
	wire [3:0] _T_171 = (muxStateEarly_6 ? out_1_6_d_bits_size : 4'h0);
	wire [3:0] _T_172 = (muxStateEarly_7 ? out_1_7_d_bits_size : 4'h0);
	wire [3:0] _T_173 = (muxStateEarly_8 ? out_1_8_d_bits_size : 4'h0);
	wire [3:0] _T_174 = _T_165 | _T_166;
	wire [3:0] _T_175 = _T_174 | _T_167;
	wire [3:0] _T_176 = _T_175 | _T_168;
	wire [3:0] _T_177 = _T_176 | _T_169;
	wire [3:0] _T_178 = _T_177 | _T_170;
	wire [3:0] _T_179 = _T_178 | _T_171;
	wire [3:0] _T_180 = _T_179 | _T_172;
	wire [1:0] _T_182 = (muxStateEarly_0 ? auto_out_0_d_bits_param : 2'h0);
	wire [1:0] _T_183 = (muxStateEarly_1 ? auto_out_1_d_bits_param : 2'h0);
	wire [1:0] _T_187 = (muxStateEarly_5 ? auto_out_5_d_bits_param : 2'h0);
	wire [1:0] _T_189 = (muxStateEarly_7 ? auto_out_7_d_bits_param : 2'h0);
	wire [1:0] _T_190 = (muxStateEarly_8 ? auto_out_8_d_bits_param : 2'h0);
	wire [1:0] _T_191 = _T_182 | _T_183;
	wire [1:0] _T_195 = _T_191 | _T_187;
	wire [1:0] _T_197 = _T_195 | _T_189;
	wire [2:0] _T_199 = (muxStateEarly_0 ? auto_out_0_d_bits_opcode : 3'h0);
	wire [2:0] _T_200 = (muxStateEarly_1 ? auto_out_1_d_bits_opcode : 3'h0);
	wire [2:0] _T_201 = (muxStateEarly_2 ? auto_out_2_d_bits_opcode : 3'h0);
	wire [2:0] _T_202 = (muxStateEarly_3 ? auto_out_3_d_bits_opcode : 3'h0);
	wire [2:0] _T_203 = (muxStateEarly_4 ? auto_out_4_d_bits_opcode : 3'h0);
	wire [2:0] _T_204 = (muxStateEarly_5 ? auto_out_5_d_bits_opcode : 3'h0);
	wire [2:0] _T_205 = (muxStateEarly_6 ? 3'h1 : 3'h0);
	wire [2:0] _T_206 = (muxStateEarly_7 ? auto_out_7_d_bits_opcode : 3'h0);
	wire [2:0] _T_207 = (muxStateEarly_8 ? auto_out_8_d_bits_opcode : 3'h0);
	wire [2:0] _T_208 = _T_199 | _T_200;
	wire [2:0] _T_209 = _T_208 | _T_201;
	wire [2:0] _T_210 = _T_209 | _T_202;
	wire [2:0] _T_211 = _T_210 | _T_203;
	wire [2:0] _T_212 = _T_211 | _T_204;
	wire [2:0] _T_213 = _T_212 | _T_205;
	wire [2:0] _T_214 = _T_213 | _T_206;
	TLMonitor_18 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	assign auto_in_a_ready = ((((((((requestAIO_0_0 & auto_out_0_a_ready) | (requestAIO_0_1 & auto_out_1_a_ready)) | (requestAIO_0_2 & auto_out_2_a_ready)) | (requestAIO_0_3 & auto_out_3_a_ready)) | (requestAIO_0_4 & auto_out_4_a_ready)) | (requestAIO_0_5 & auto_out_5_a_ready)) | (requestAIO_0_6 & auto_out_6_a_ready)) | (requestAIO_0_7 & auto_out_7_a_ready)) | (requestAIO_0_8 & auto_out_8_a_ready);
	assign auto_in_d_valid = (idle ? _T_45 : _sink_ACancel_earlyValid_T_24);
	assign auto_in_d_bits_opcode = _T_214 | _T_207;
	assign auto_in_d_bits_param = _T_197 | _T_190;
	assign auto_in_d_bits_size = _T_180 | _T_173;
	assign auto_in_d_bits_source = _T_163 | _T_156;
	assign auto_in_d_bits_sink = ((((muxStateEarly_0 & auto_out_0_d_bits_sink) | (muxStateEarly_1 & auto_out_1_d_bits_sink)) | (muxStateEarly_5 & auto_out_5_d_bits_sink)) | (muxStateEarly_7 & auto_out_7_d_bits_sink)) | (muxStateEarly_8 & auto_out_8_d_bits_sink);
	assign auto_in_d_bits_denied = ((((muxStateEarly_0 & auto_out_0_d_bits_denied) | (muxStateEarly_1 & auto_out_1_d_bits_denied)) | (muxStateEarly_5 & auto_out_5_d_bits_denied)) | (muxStateEarly_7 & auto_out_7_d_bits_denied)) | (muxStateEarly_8 & auto_out_8_d_bits_denied);
	assign auto_in_d_bits_data = _T_112 | _T_105;
	assign auto_in_d_bits_corrupt = ((((muxStateEarly_0 & auto_out_0_d_bits_corrupt) | (muxStateEarly_1 & auto_out_1_d_bits_corrupt)) | (muxStateEarly_5 & auto_out_5_d_bits_corrupt)) | (muxStateEarly_7 & auto_out_7_d_bits_corrupt)) | (muxStateEarly_8 & auto_out_8_d_bits_corrupt);
	assign auto_out_8_a_valid = auto_in_a_valid & requestAIO_0_8;
	assign auto_out_8_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_8_a_bits_param = auto_in_a_bits_param;
	assign auto_out_8_a_bits_size = auto_in_a_bits_size[2:0];
	assign auto_out_8_a_bits_source = auto_in_a_bits_source;
	assign auto_out_8_a_bits_address = auto_in_a_bits_address[20:0];
	assign auto_out_8_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_8_a_bits_data = auto_in_a_bits_data;
	assign auto_out_8_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_8_d_ready = auto_in_d_ready & allowed_8;
	assign auto_out_7_a_valid = auto_in_a_valid & requestAIO_0_7;
	assign auto_out_7_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_7_a_bits_param = auto_in_a_bits_param;
	assign auto_out_7_a_bits_size = auto_in_a_bits_size[2:0];
	assign auto_out_7_a_bits_source = auto_in_a_bits_source;
	assign auto_out_7_a_bits_address = auto_in_a_bits_address[20:0];
	assign auto_out_7_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_7_a_bits_data = auto_in_a_bits_data;
	assign auto_out_7_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_7_d_ready = auto_in_d_ready & allowed_7;
	assign auto_out_6_a_valid = auto_in_a_valid & requestAIO_0_6;
	assign auto_out_6_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_6_a_bits_param = auto_in_a_bits_param;
	assign auto_out_6_a_bits_size = auto_in_a_bits_size[2:0];
	assign auto_out_6_a_bits_source = auto_in_a_bits_source;
	assign auto_out_6_a_bits_address = auto_in_a_bits_address[16:0];
	assign auto_out_6_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_6_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_6_d_ready = auto_in_d_ready & allowed_6;
	assign auto_out_5_a_valid = auto_in_a_valid & requestAIO_0_5;
	assign auto_out_5_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_5_a_bits_param = auto_in_a_bits_param;
	assign auto_out_5_a_bits_size = auto_in_a_bits_size[2:0];
	assign auto_out_5_a_bits_source = auto_in_a_bits_source;
	assign auto_out_5_a_bits_address = auto_in_a_bits_address;
	assign auto_out_5_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_5_a_bits_data = auto_in_a_bits_data;
	assign auto_out_5_d_ready = auto_in_d_ready & allowed_5;
	assign auto_out_4_a_valid = auto_in_a_valid & requestAIO_0_4;
	assign auto_out_4_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_4_a_bits_param = auto_in_a_bits_param;
	assign auto_out_4_a_bits_size = auto_in_a_bits_size[2:0];
	assign auto_out_4_a_bits_source = auto_in_a_bits_source;
	assign auto_out_4_a_bits_address = auto_in_a_bits_address[11:0];
	assign auto_out_4_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_4_a_bits_data = auto_in_a_bits_data;
	assign auto_out_4_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_4_d_ready = auto_in_d_ready & allowed_4;
	assign auto_out_3_a_valid = auto_in_a_valid & requestAIO_0_3;
	assign auto_out_3_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_3_a_bits_param = auto_in_a_bits_param;
	assign auto_out_3_a_bits_size = auto_in_a_bits_size[2:0];
	assign auto_out_3_a_bits_source = auto_in_a_bits_source;
	assign auto_out_3_a_bits_address = auto_in_a_bits_address[25:0];
	assign auto_out_3_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_3_a_bits_data = auto_in_a_bits_data;
	assign auto_out_3_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_3_d_ready = auto_in_d_ready & allowed_3;
	assign auto_out_2_a_valid = auto_in_a_valid & requestAIO_0_2;
	assign auto_out_2_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_2_a_bits_param = auto_in_a_bits_param;
	assign auto_out_2_a_bits_size = auto_in_a_bits_size[2:0];
	assign auto_out_2_a_bits_source = auto_in_a_bits_source;
	assign auto_out_2_a_bits_address = auto_in_a_bits_address[27:0];
	assign auto_out_2_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_2_a_bits_data = auto_in_a_bits_data;
	assign auto_out_2_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_2_d_ready = auto_in_d_ready & allowed_2;
	assign auto_out_1_a_valid = auto_in_a_valid & requestAIO_0_1;
	assign auto_out_1_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_1_a_bits_param = auto_in_a_bits_param;
	assign auto_out_1_a_bits_size = auto_in_a_bits_size[2:0];
	assign auto_out_1_a_bits_source = auto_in_a_bits_source;
	assign auto_out_1_a_bits_address = auto_in_a_bits_address[30:0];
	assign auto_out_1_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_1_a_bits_data = auto_in_a_bits_data;
	assign auto_out_1_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_1_d_ready = auto_in_d_ready & allowed_1;
	assign auto_out_0_a_valid = auto_in_a_valid & requestAIO_0_0;
	assign auto_out_0_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_0_a_bits_param = auto_in_a_bits_param;
	assign auto_out_0_a_bits_size = auto_in_a_bits_size;
	assign auto_out_0_a_bits_source = auto_in_a_bits_source;
	assign auto_out_0_a_bits_address = auto_in_a_bits_address[13:0];
	assign auto_out_0_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_0_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_0_d_ready = auto_in_d_ready & allowed_0;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = ((((((((requestAIO_0_0 & auto_out_0_a_ready) | (requestAIO_0_1 & auto_out_1_a_ready)) | (requestAIO_0_2 & auto_out_2_a_ready)) | (requestAIO_0_3 & auto_out_3_a_ready)) | (requestAIO_0_4 & auto_out_4_a_ready)) | (requestAIO_0_5 & auto_out_5_a_ready)) | (requestAIO_0_6 & auto_out_6_a_ready)) | (requestAIO_0_7 & auto_out_7_a_ready)) | (requestAIO_0_8 & auto_out_8_a_ready);
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = (idle ? _T_45 : _sink_ACancel_earlyValid_T_24);
	assign monitor_io_in_d_bits_opcode = _T_214 | _T_207;
	assign monitor_io_in_d_bits_param = _T_197 | _T_190;
	assign monitor_io_in_d_bits_size = _T_180 | _T_173;
	assign monitor_io_in_d_bits_source = _T_163 | _T_156;
	assign monitor_io_in_d_bits_sink = ((((muxStateEarly_0 & auto_out_0_d_bits_sink) | (muxStateEarly_1 & auto_out_1_d_bits_sink)) | (muxStateEarly_5 & auto_out_5_d_bits_sink)) | (muxStateEarly_7 & auto_out_7_d_bits_sink)) | (muxStateEarly_8 & auto_out_8_d_bits_sink);
	assign monitor_io_in_d_bits_denied = ((((muxStateEarly_0 & auto_out_0_d_bits_denied) | (muxStateEarly_1 & auto_out_1_d_bits_denied)) | (muxStateEarly_5 & auto_out_5_d_bits_denied)) | (muxStateEarly_7 & auto_out_7_d_bits_denied)) | (muxStateEarly_8 & auto_out_8_d_bits_denied);
	assign monitor_io_in_d_bits_corrupt = ((((muxStateEarly_0 & auto_out_0_d_bits_corrupt) | (muxStateEarly_1 & auto_out_1_d_bits_corrupt)) | (muxStateEarly_5 & auto_out_5_d_bits_corrupt)) | (muxStateEarly_7 & auto_out_7_d_bits_corrupt)) | (muxStateEarly_8 & auto_out_8_d_bits_corrupt);
	always @(posedge clock) begin
		if (reset)
			beatsLeft <= 10'h000;
		else if (latch)
			beatsLeft <= initBeats;
		else
			beatsLeft <= _beatsLeft_T_4;
		if (reset)
			readys_mask <= 9'h1ff;
		else if (latch & |readys_valid)
			readys_mask <= _readys_mask_T_12;
		if (reset)
			state_0 <= 1'h0;
		else if (idle)
			state_0 <= earlyWinner_0;
		if (reset)
			state_1 <= 1'h0;
		else if (idle)
			state_1 <= earlyWinner_1;
		if (reset)
			state_2 <= 1'h0;
		else if (idle)
			state_2 <= earlyWinner_2;
		if (reset)
			state_3 <= 1'h0;
		else if (idle)
			state_3 <= earlyWinner_3;
		if (reset)
			state_4 <= 1'h0;
		else if (idle)
			state_4 <= earlyWinner_4;
		if (reset)
			state_5 <= 1'h0;
		else if (idle)
			state_5 <= earlyWinner_5;
		if (reset)
			state_6 <= 1'h0;
		else if (idle)
			state_6 <= earlyWinner_6;
		if (reset)
			state_7 <= 1'h0;
		else if (idle)
			state_7 <= earlyWinner_7;
		if (reset)
			state_8 <= 1'h0;
		else if (idle)
			state_8 <= earlyWinner_8;
	end
endmodule
module TLMonitor_19 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire _T_44 = io_in_a_bits_size <= 4'hc;
	wire _T_53 = _T_44 & source_ok;
	wire [32:0] _T_59 = $signed(_T_7) & -33'sh000005000;
	wire _T_60 = $signed(_T_59) == 33'sh000000000;
	wire [31:0] _T_61 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_62 = {1'b0, $signed(_T_61)};
	wire [32:0] _T_64 = $signed(_T_62) & -33'sh000001000;
	wire _T_65 = $signed(_T_64) == 33'sh000000000;
	wire [31:0] _T_66 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_67 = {1'b0, $signed(_T_66)};
	wire [32:0] _T_69 = $signed(_T_67) & -33'sh000010000;
	wire _T_70 = $signed(_T_69) == 33'sh000000000;
	wire [31:0] _T_71 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_72 = {1'b0, $signed(_T_71)};
	wire [32:0] _T_74 = $signed(_T_72) & -33'sh000010000;
	wire _T_75 = $signed(_T_74) == 33'sh000000000;
	wire [31:0] _T_76 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_77 = {1'b0, $signed(_T_76)};
	wire [32:0] _T_79 = $signed(_T_77) & -33'sh000011000;
	wire _T_80 = $signed(_T_79) == 33'sh000000000;
	wire [31:0] _T_81 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_82 = {1'b0, $signed(_T_81)};
	wire [32:0] _T_84 = $signed(_T_82) & -33'sh000010000;
	wire _T_85 = $signed(_T_84) == 33'sh000000000;
	wire [31:0] _T_86 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_87 = {1'b0, $signed(_T_86)};
	wire [32:0] _T_89 = $signed(_T_87) & -33'sh004000000;
	wire _T_90 = $signed(_T_89) == 33'sh000000000;
	wire [31:0] _T_91 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_92 = {1'b0, $signed(_T_91)};
	wire [32:0] _T_94 = $signed(_T_92) & -33'sh000001000;
	wire _T_95 = $signed(_T_94) == 33'sh000000000;
	wire [31:0] _T_96 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_97 = {1'b0, $signed(_T_96)};
	wire [32:0] _T_99 = $signed(_T_97) & -33'sh000001000;
	wire _T_100 = $signed(_T_99) == 33'sh000000000;
	wire [31:0] _T_101 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_102 = {1'b0, $signed(_T_101)};
	wire [32:0] _T_104 = $signed(_T_102) & -33'sh000004000;
	wire _T_105 = $signed(_T_104) == 33'sh000000000;
	wire _T_200 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_204 = ~io_in_a_bits_mask;
	wire _T_205 = _T_204 == 4'h0;
	wire _T_209 = ~io_in_a_bits_corrupt;
	wire _T_213 = io_in_a_bits_opcode == 3'h7;
	wire _T_375 = io_in_a_bits_param != 3'h0;
	wire _T_388 = io_in_a_bits_opcode == 3'h4;
	wire _T_413 = _T_44 & _T_65;
	wire _T_415 = io_in_a_bits_size <= 4'h6;
	wire _T_470 = (((((((_T_60 | _T_70) | _T_75) | _T_80) | _T_85) | _T_90) | _T_95) | _T_100) | _T_105;
	wire _T_471 = _T_415 & _T_470;
	wire _T_473 = _T_413 | _T_471;
	wire _T_483 = io_in_a_bits_param == 3'h0;
	wire _T_487 = io_in_a_bits_mask == mask;
	wire _T_495 = io_in_a_bits_opcode == 3'h0;
	wire _T_562 = (((((_T_60 | _T_80) | _T_85) | _T_90) | _T_95) | _T_100) | _T_105;
	wire _T_563 = _T_415 & _T_562;
	wire _T_578 = _T_413 | _T_563;
	wire _T_580 = _T_53 & _T_578;
	wire _T_598 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_697 = ~mask;
	wire [3:0] _T_698 = io_in_a_bits_mask & _T_697;
	wire _T_699 = _T_698 == 4'h0;
	wire _T_703 = io_in_a_bits_opcode == 3'h2;
	wire _T_717 = io_in_a_bits_size <= 4'h2;
	wire [31:0] _T_725 = io_in_a_bits_address ^ 32'h00004000;
	wire [32:0] _T_726 = {1'b0, $signed(_T_725)};
	wire [32:0] _T_728 = $signed(_T_726) & -33'sh000001000;
	wire _T_729 = $signed(_T_728) == 33'sh000000000;
	wire _T_742 = ((_T_65 | _T_729) | _T_95) | _T_100;
	wire _T_743 = _T_717 & _T_742;
	wire _T_781 = 4'h2 == io_in_a_bits_size;
	wire _T_788 = _T_781 & _T_105;
	wire _T_791 = _T_743 | _T_788;
	wire _T_792 = _T_53 & _T_791;
	wire _T_802 = io_in_a_bits_param <= 3'h4;
	wire _T_810 = io_in_a_bits_opcode == 3'h3;
	wire _T_909 = io_in_a_bits_param <= 3'h3;
	wire _T_917 = io_in_a_bits_opcode == 3'h5;
	wire _T_997 = _T_53 & _T_413;
	wire _T_1007 = io_in_a_bits_param <= 3'h1;
	wire _T_1019 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_1023 = io_in_d_bits_opcode == 3'h6;
	wire _T_1027 = io_in_d_bits_size >= 4'h2;
	wire _T_1031 = io_in_d_bits_param == 2'h0;
	wire _T_1035 = ~io_in_d_bits_corrupt;
	wire _T_1039 = ~io_in_d_bits_denied;
	wire _T_1043 = io_in_d_bits_opcode == 3'h4;
	wire _T_1054 = io_in_d_bits_param <= 2'h2;
	wire _T_1058 = io_in_d_bits_param != 2'h2;
	wire _T_1071 = io_in_d_bits_opcode == 3'h5;
	wire _T_1091 = _T_1039 | io_in_d_bits_corrupt;
	wire _T_1100 = io_in_d_bits_opcode == 3'h0;
	wire _T_1117 = io_in_d_bits_opcode == 3'h1;
	wire _T_1135 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg [2:0] source;
	reg [31:0] address;
	wire _T_1165 = io_in_a_valid & ~a_first;
	wire _T_1166 = io_in_a_bits_opcode == opcode;
	wire _T_1170 = io_in_a_bits_param == param;
	wire _T_1174 = io_in_a_bits_size == size;
	wire _T_1178 = io_in_a_bits_source == source;
	wire _T_1182 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_1189 = io_in_d_valid & ~d_first;
	wire _T_1190 = io_in_d_bits_opcode == opcode_1;
	wire _T_1194 = io_in_d_bits_param == param_1;
	wire _T_1198 = io_in_d_bits_size == size_1;
	wire _T_1202 = io_in_d_bits_source == source_1;
	wire _T_1206 = io_in_d_bits_sink == sink;
	wire _T_1210 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [39:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [5:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0};
	wire [39:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T;
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [39:0] _GEN_75 = {24'd0, _a_size_lookup_T_5};
	wire [39:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_75;
	wire [39:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[39:1]};
	wire _T_1216 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire [7:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire _T_1219 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [4:0] _GEN_77 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_77};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [5:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [67:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [67:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire [4:0] _T_1221 = inflight >> io_in_a_bits_source;
	wire _T_1223 = ~_T_1221[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [67:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 68'h00000000000000000);
	wire _T_1227 = io_in_d_valid & d_first_1;
	wire _T_1229 = ~_T_1023;
	wire _T_1230 = (io_in_d_valid & d_first_1) & ~_T_1023;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [7:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_1023 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [78:0] _GEN_4 = {63'd0, _a_size_lookup_T_5};
	wire [78:0] _d_sizes_clr_T_5 = _GEN_4 << _a_size_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_1229 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1229 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [78:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1229 ? _d_sizes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_1216 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_1240 = inflight >> io_in_d_bits_source;
	wire _T_1242 = _T_1240[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1247 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1248 = (io_in_d_bits_opcode == _GEN_32) | _T_1247;
	wire _T_1252 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1259 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1260 = (io_in_d_bits_opcode == _GEN_48) | _T_1259;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_79 = {4'd0, io_in_d_bits_size};
	wire _T_1264 = _GEN_79 == a_size_lookup;
	wire _T_1274 = (((_T_1227 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_1229;
	wire _T_1276 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set_wo_ready = _GEN_15[4:0];
	wire [4:0] d_clr_wo_ready = _GEN_21[4:0];
	wire _T_1283 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [39:0] a_sizes_set = _GEN_20[39:0];
	wire [39:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [39:0] d_sizes_clr = _GEN_24[39:0];
	wire [39:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [39:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1292 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [39:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [39:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T;
	wire [39:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_75;
	wire [39:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[39:1]};
	wire _T_1318 = (io_in_d_valid & d_first_2) & _T_1023;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_1023 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_1023 ? _d_sizes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_1326 = inflight_1 >> io_in_d_bits_source;
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1336 = _GEN_79 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [39:0] d_sizes_clr_1 = _GEN_69[39:0];
	wire [39:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [39:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	reg [31:0] watchdog_1;
	wire _T_1361 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 40'h0000000000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 40'h0000000000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Queue_8 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_data,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [3:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [31:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input [31:0] io_enq_bits_data;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [3:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [31:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire [31:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg [2:0] ram_opcode [0:1];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [2:0] ram_param [0:1];
	wire ram_param_io_deq_bits_MPORT_en;
	wire ram_param_io_deq_bits_MPORT_addr;
	wire [2:0] ram_param_io_deq_bits_MPORT_data;
	wire [2:0] ram_param_MPORT_data;
	wire ram_param_MPORT_addr;
	wire ram_param_MPORT_mask;
	wire ram_param_MPORT_en;
	reg [3:0] ram_size [0:1];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [3:0] ram_size_io_deq_bits_MPORT_data;
	wire [3:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg [2:0] ram_source [0:1];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire [2:0] ram_source_io_deq_bits_MPORT_data;
	wire [2:0] ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg [31:0] ram_address [0:1];
	wire ram_address_io_deq_bits_MPORT_en;
	wire ram_address_io_deq_bits_MPORT_addr;
	wire [31:0] ram_address_io_deq_bits_MPORT_data;
	wire [31:0] ram_address_MPORT_data;
	wire ram_address_MPORT_addr;
	wire ram_address_MPORT_mask;
	wire ram_address_MPORT_en;
	reg [3:0] ram_mask [0:1];
	wire ram_mask_io_deq_bits_MPORT_en;
	wire ram_mask_io_deq_bits_MPORT_addr;
	wire [3:0] ram_mask_io_deq_bits_MPORT_data;
	wire [3:0] ram_mask_MPORT_data;
	wire ram_mask_MPORT_addr;
	wire ram_mask_MPORT_mask;
	wire ram_mask_MPORT_en;
	reg [31:0] ram_data [0:1];
	wire ram_data_io_deq_bits_MPORT_en;
	wire ram_data_io_deq_bits_MPORT_addr;
	wire [31:0] ram_data_io_deq_bits_MPORT_data;
	wire [31:0] ram_data_MPORT_data;
	wire ram_data_MPORT_addr;
	wire ram_data_MPORT_mask;
	wire ram_data_MPORT_en;
	reg ram_corrupt [0:1];
	wire ram_corrupt_io_deq_bits_MPORT_en;
	wire ram_corrupt_io_deq_bits_MPORT_addr;
	wire ram_corrupt_io_deq_bits_MPORT_data;
	wire ram_corrupt_MPORT_data;
	wire ram_corrupt_MPORT_addr;
	wire ram_corrupt_MPORT_mask;
	wire ram_corrupt_MPORT_en;
	reg value;
	reg value_1;
	reg maybe_full;
	wire ptr_match = value == value_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = value;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_param_io_deq_bits_MPORT_en = 1'h1;
	assign ram_param_io_deq_bits_MPORT_addr = value_1;
	assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr];
	assign ram_param_MPORT_data = io_enq_bits_param;
	assign ram_param_MPORT_addr = value;
	assign ram_param_MPORT_mask = 1'h1;
	assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = value_1;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = value;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = value_1;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = value;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_address_io_deq_bits_MPORT_en = 1'h1;
	assign ram_address_io_deq_bits_MPORT_addr = value_1;
	assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr];
	assign ram_address_MPORT_data = io_enq_bits_address;
	assign ram_address_MPORT_addr = value;
	assign ram_address_MPORT_mask = 1'h1;
	assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
	assign ram_mask_io_deq_bits_MPORT_addr = value_1;
	assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr];
	assign ram_mask_MPORT_data = io_enq_bits_mask;
	assign ram_mask_MPORT_addr = value;
	assign ram_mask_MPORT_mask = 1'h1;
	assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_data_io_deq_bits_MPORT_en = 1'h1;
	assign ram_data_io_deq_bits_MPORT_addr = value_1;
	assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr];
	assign ram_data_MPORT_data = io_enq_bits_data;
	assign ram_data_MPORT_addr = value;
	assign ram_data_MPORT_mask = 1'h1;
	assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
	assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
	assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr];
	assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
	assign ram_corrupt_MPORT_addr = value;
	assign ram_corrupt_MPORT_mask = 1'h1;
	assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data;
	assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data;
	assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data;
	assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_param_MPORT_en & ram_param_MPORT_mask)
			ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (ram_address_MPORT_en & ram_address_MPORT_mask)
			ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data;
		if (ram_mask_MPORT_en & ram_mask_MPORT_mask)
			ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data;
		if (ram_data_MPORT_en & ram_data_MPORT_mask)
			ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data;
		if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask)
			ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data;
		if (reset)
			value <= 1'h0;
		else if (do_enq)
			value <= value + 1'h1;
		if (reset)
			value_1 <= 1'h0;
		else if (do_deq)
			value_1 <= value_1 + 1'h1;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module Queue_9 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_sink,
	io_enq_bits_denied,
	io_enq_bits_data,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_sink,
	io_deq_bits_denied,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [1:0] io_enq_bits_param;
	input [3:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input io_enq_bits_sink;
	input io_enq_bits_denied;
	input [31:0] io_enq_bits_data;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [1:0] io_deq_bits_param;
	output wire [3:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire io_deq_bits_sink;
	output wire io_deq_bits_denied;
	output wire [31:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg [2:0] ram_opcode [0:1];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [1:0] ram_param [0:1];
	wire ram_param_io_deq_bits_MPORT_en;
	wire ram_param_io_deq_bits_MPORT_addr;
	wire [1:0] ram_param_io_deq_bits_MPORT_data;
	wire [1:0] ram_param_MPORT_data;
	wire ram_param_MPORT_addr;
	wire ram_param_MPORT_mask;
	wire ram_param_MPORT_en;
	reg [3:0] ram_size [0:1];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [3:0] ram_size_io_deq_bits_MPORT_data;
	wire [3:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg [2:0] ram_source [0:1];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire [2:0] ram_source_io_deq_bits_MPORT_data;
	wire [2:0] ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg ram_sink [0:1];
	wire ram_sink_io_deq_bits_MPORT_en;
	wire ram_sink_io_deq_bits_MPORT_addr;
	wire ram_sink_io_deq_bits_MPORT_data;
	wire ram_sink_MPORT_data;
	wire ram_sink_MPORT_addr;
	wire ram_sink_MPORT_mask;
	wire ram_sink_MPORT_en;
	reg ram_denied [0:1];
	wire ram_denied_io_deq_bits_MPORT_en;
	wire ram_denied_io_deq_bits_MPORT_addr;
	wire ram_denied_io_deq_bits_MPORT_data;
	wire ram_denied_MPORT_data;
	wire ram_denied_MPORT_addr;
	wire ram_denied_MPORT_mask;
	wire ram_denied_MPORT_en;
	reg [31:0] ram_data [0:1];
	wire ram_data_io_deq_bits_MPORT_en;
	wire ram_data_io_deq_bits_MPORT_addr;
	wire [31:0] ram_data_io_deq_bits_MPORT_data;
	wire [31:0] ram_data_MPORT_data;
	wire ram_data_MPORT_addr;
	wire ram_data_MPORT_mask;
	wire ram_data_MPORT_en;
	reg ram_corrupt [0:1];
	wire ram_corrupt_io_deq_bits_MPORT_en;
	wire ram_corrupt_io_deq_bits_MPORT_addr;
	wire ram_corrupt_io_deq_bits_MPORT_data;
	wire ram_corrupt_MPORT_data;
	wire ram_corrupt_MPORT_addr;
	wire ram_corrupt_MPORT_mask;
	wire ram_corrupt_MPORT_en;
	reg value;
	reg value_1;
	reg maybe_full;
	wire ptr_match = value == value_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = value;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_param_io_deq_bits_MPORT_en = 1'h1;
	assign ram_param_io_deq_bits_MPORT_addr = value_1;
	assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr];
	assign ram_param_MPORT_data = io_enq_bits_param;
	assign ram_param_MPORT_addr = value;
	assign ram_param_MPORT_mask = 1'h1;
	assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = value_1;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = value;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = value_1;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = value;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_sink_io_deq_bits_MPORT_en = 1'h1;
	assign ram_sink_io_deq_bits_MPORT_addr = value_1;
	assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr];
	assign ram_sink_MPORT_data = io_enq_bits_sink;
	assign ram_sink_MPORT_addr = value;
	assign ram_sink_MPORT_mask = 1'h1;
	assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_denied_io_deq_bits_MPORT_en = 1'h1;
	assign ram_denied_io_deq_bits_MPORT_addr = value_1;
	assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr];
	assign ram_denied_MPORT_data = io_enq_bits_denied;
	assign ram_denied_MPORT_addr = value;
	assign ram_denied_MPORT_mask = 1'h1;
	assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_data_io_deq_bits_MPORT_en = 1'h1;
	assign ram_data_io_deq_bits_MPORT_addr = value_1;
	assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr];
	assign ram_data_MPORT_data = io_enq_bits_data;
	assign ram_data_MPORT_addr = value;
	assign ram_data_MPORT_mask = 1'h1;
	assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
	assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
	assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr];
	assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
	assign ram_corrupt_MPORT_addr = value;
	assign ram_corrupt_MPORT_mask = 1'h1;
	assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data;
	assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data;
	assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data;
	assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_param_MPORT_en & ram_param_MPORT_mask)
			ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (ram_sink_MPORT_en & ram_sink_MPORT_mask)
			ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data;
		if (ram_denied_MPORT_en & ram_denied_MPORT_mask)
			ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data;
		if (ram_data_MPORT_en & ram_data_MPORT_mask)
			ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data;
		if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask)
			ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data;
		if (reset)
			value <= 1'h0;
		else if (do_enq)
			value <= value + 1'h1;
		if (reset)
			value_1 <= 1'h0;
		else if (do_deq)
			value_1 <= value_1 + 1'h1;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module TLBuffer_6 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [31:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [3:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire bundleOut_0_a_q_clock;
	wire bundleOut_0_a_q_reset;
	wire bundleOut_0_a_q_io_enq_ready;
	wire bundleOut_0_a_q_io_enq_valid;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_param;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_size;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_source;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_data;
	wire bundleOut_0_a_q_io_enq_bits_corrupt;
	wire bundleOut_0_a_q_io_deq_ready;
	wire bundleOut_0_a_q_io_deq_valid;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_param;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_size;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_source;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_data;
	wire bundleOut_0_a_q_io_deq_bits_corrupt;
	wire bundleIn_0_d_q_clock;
	wire bundleIn_0_d_q_reset;
	wire bundleIn_0_d_q_io_enq_ready;
	wire bundleIn_0_d_q_io_enq_valid;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_enq_bits_param;
	wire [3:0] bundleIn_0_d_q_io_enq_bits_size;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_source;
	wire bundleIn_0_d_q_io_enq_bits_sink;
	wire bundleIn_0_d_q_io_enq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_enq_bits_data;
	wire bundleIn_0_d_q_io_enq_bits_corrupt;
	wire bundleIn_0_d_q_io_deq_ready;
	wire bundleIn_0_d_q_io_deq_valid;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_param;
	wire [3:0] bundleIn_0_d_q_io_deq_bits_size;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_source;
	wire bundleIn_0_d_q_io_deq_bits_sink;
	wire bundleIn_0_d_q_io_deq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_deq_bits_data;
	wire bundleIn_0_d_q_io_deq_bits_corrupt;
	TLMonitor_19 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Queue_8 bundleOut_0_a_q(
		.clock(bundleOut_0_a_q_clock),
		.reset(bundleOut_0_a_q_reset),
		.io_enq_ready(bundleOut_0_a_q_io_enq_ready),
		.io_enq_valid(bundleOut_0_a_q_io_enq_valid),
		.io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
		.io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
		.io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
		.io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
		.io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
		.io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleOut_0_a_q_io_deq_ready),
		.io_deq_valid(bundleOut_0_a_q_io_deq_valid),
		.io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
		.io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
		.io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
		.io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
		.io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
		.io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
	);
	Queue_9 bundleIn_0_d_q(
		.clock(bundleIn_0_d_q_clock),
		.reset(bundleIn_0_d_q_reset),
		.io_enq_ready(bundleIn_0_d_q_io_enq_ready),
		.io_enq_valid(bundleIn_0_d_q_io_enq_valid),
		.io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
		.io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
		.io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
		.io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
		.io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
		.io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleIn_0_d_q_io_deq_ready),
		.io_deq_valid(bundleIn_0_d_q_io_deq_valid),
		.io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
		.io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
		.io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
		.io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
		.io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
		.io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data;
	assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid;
	assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode;
	assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param;
	assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size;
	assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source;
	assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address;
	assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask;
	assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data;
	assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt;
	assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign bundleOut_0_a_q_clock = clock;
	assign bundleOut_0_a_q_reset = reset;
	assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid;
	assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param;
	assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size;
	assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source;
	assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address;
	assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask;
	assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data;
	assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready;
	assign bundleIn_0_d_q_clock = clock;
	assign bundleIn_0_d_q_reset = reset;
	assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid;
	assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign bundleIn_0_d_q_io_enq_bits_param = auto_out_d_bits_param;
	assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size;
	assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source;
	assign bundleIn_0_d_q_io_enq_bits_sink = auto_out_d_bits_sink;
	assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied;
	assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data;
	assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt;
	assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready;
endmodule
module TLMonitor_20 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire _T_44 = io_in_a_bits_size <= 4'hc;
	wire _T_53 = _T_44 & source_ok;
	wire [32:0] _T_59 = $signed(_T_7) & -33'sh000005000;
	wire _T_60 = $signed(_T_59) == 33'sh000000000;
	wire [31:0] _T_61 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_62 = {1'b0, $signed(_T_61)};
	wire [32:0] _T_64 = $signed(_T_62) & -33'sh000001000;
	wire _T_65 = $signed(_T_64) == 33'sh000000000;
	wire [31:0] _T_66 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_67 = {1'b0, $signed(_T_66)};
	wire [32:0] _T_69 = $signed(_T_67) & -33'sh000010000;
	wire _T_70 = $signed(_T_69) == 33'sh000000000;
	wire [31:0] _T_71 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_72 = {1'b0, $signed(_T_71)};
	wire [32:0] _T_74 = $signed(_T_72) & -33'sh000010000;
	wire _T_75 = $signed(_T_74) == 33'sh000000000;
	wire [31:0] _T_76 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_77 = {1'b0, $signed(_T_76)};
	wire [32:0] _T_79 = $signed(_T_77) & -33'sh000011000;
	wire _T_80 = $signed(_T_79) == 33'sh000000000;
	wire [31:0] _T_81 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_82 = {1'b0, $signed(_T_81)};
	wire [32:0] _T_84 = $signed(_T_82) & -33'sh000010000;
	wire _T_85 = $signed(_T_84) == 33'sh000000000;
	wire [31:0] _T_86 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_87 = {1'b0, $signed(_T_86)};
	wire [32:0] _T_89 = $signed(_T_87) & -33'sh004000000;
	wire _T_90 = $signed(_T_89) == 33'sh000000000;
	wire [31:0] _T_91 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_92 = {1'b0, $signed(_T_91)};
	wire [32:0] _T_94 = $signed(_T_92) & -33'sh000001000;
	wire _T_95 = $signed(_T_94) == 33'sh000000000;
	wire [31:0] _T_96 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_97 = {1'b0, $signed(_T_96)};
	wire [32:0] _T_99 = $signed(_T_97) & -33'sh000001000;
	wire _T_100 = $signed(_T_99) == 33'sh000000000;
	wire [31:0] _T_101 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_102 = {1'b0, $signed(_T_101)};
	wire [32:0] _T_104 = $signed(_T_102) & -33'sh000004000;
	wire _T_105 = $signed(_T_104) == 33'sh000000000;
	wire _T_200 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_204 = ~io_in_a_bits_mask;
	wire _T_205 = _T_204 == 4'h0;
	wire _T_209 = ~io_in_a_bits_corrupt;
	wire _T_213 = io_in_a_bits_opcode == 3'h7;
	wire _T_375 = io_in_a_bits_param != 3'h0;
	wire _T_388 = io_in_a_bits_opcode == 3'h4;
	wire _T_413 = _T_44 & _T_65;
	wire _T_415 = io_in_a_bits_size <= 4'h6;
	wire _T_470 = (((((((_T_60 | _T_70) | _T_75) | _T_80) | _T_85) | _T_90) | _T_95) | _T_100) | _T_105;
	wire _T_471 = _T_415 & _T_470;
	wire _T_473 = _T_413 | _T_471;
	wire _T_483 = io_in_a_bits_param == 3'h0;
	wire _T_487 = io_in_a_bits_mask == mask;
	wire _T_495 = io_in_a_bits_opcode == 3'h0;
	wire _T_562 = (((((_T_60 | _T_80) | _T_85) | _T_90) | _T_95) | _T_100) | _T_105;
	wire _T_563 = _T_415 & _T_562;
	wire _T_578 = _T_413 | _T_563;
	wire _T_580 = _T_53 & _T_578;
	wire _T_598 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_697 = ~mask;
	wire [3:0] _T_698 = io_in_a_bits_mask & _T_697;
	wire _T_699 = _T_698 == 4'h0;
	wire _T_703 = io_in_a_bits_opcode == 3'h2;
	wire _T_717 = io_in_a_bits_size <= 4'h2;
	wire _T_766 = ((((((_T_60 | _T_65) | _T_80) | _T_85) | _T_90) | _T_95) | _T_100) | _T_105;
	wire _T_767 = _T_717 & _T_766;
	wire _T_783 = _T_53 & _T_767;
	wire _T_793 = io_in_a_bits_param <= 3'h4;
	wire _T_801 = io_in_a_bits_opcode == 3'h3;
	wire _T_891 = io_in_a_bits_param <= 3'h3;
	wire _T_899 = io_in_a_bits_opcode == 3'h5;
	wire _T_979 = _T_53 & _T_413;
	wire _T_989 = io_in_a_bits_param <= 3'h1;
	wire _T_1001 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_1005 = io_in_d_bits_opcode == 3'h6;
	wire _T_1009 = io_in_d_bits_size >= 4'h2;
	wire _T_1013 = io_in_d_bits_param == 2'h0;
	wire _T_1017 = ~io_in_d_bits_corrupt;
	wire _T_1021 = ~io_in_d_bits_denied;
	wire _T_1025 = io_in_d_bits_opcode == 3'h4;
	wire _T_1036 = io_in_d_bits_param <= 2'h2;
	wire _T_1040 = io_in_d_bits_param != 2'h2;
	wire _T_1053 = io_in_d_bits_opcode == 3'h5;
	wire _T_1073 = _T_1021 | io_in_d_bits_corrupt;
	wire _T_1082 = io_in_d_bits_opcode == 3'h0;
	wire _T_1099 = io_in_d_bits_opcode == 3'h1;
	wire _T_1117 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg [2:0] source;
	reg [31:0] address;
	wire _T_1147 = io_in_a_valid & ~a_first;
	wire _T_1148 = io_in_a_bits_opcode == opcode;
	wire _T_1152 = io_in_a_bits_param == param;
	wire _T_1156 = io_in_a_bits_size == size;
	wire _T_1160 = io_in_a_bits_source == source;
	wire _T_1164 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_1171 = io_in_d_valid & ~d_first;
	wire _T_1172 = io_in_d_bits_opcode == opcode_1;
	wire _T_1176 = io_in_d_bits_param == param_1;
	wire _T_1180 = io_in_d_bits_size == size_1;
	wire _T_1184 = io_in_d_bits_source == source_1;
	wire _T_1188 = io_in_d_bits_sink == sink;
	wire _T_1192 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [39:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [5:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0};
	wire [39:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T;
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [39:0] _GEN_75 = {24'd0, _a_size_lookup_T_5};
	wire [39:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_75;
	wire [39:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[39:1]};
	wire _T_1198 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire [7:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire _T_1201 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [4:0] _GEN_77 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_77};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [5:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [67:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [67:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire [4:0] _T_1203 = inflight >> io_in_a_bits_source;
	wire _T_1205 = ~_T_1203[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [67:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 68'h00000000000000000);
	wire _T_1209 = io_in_d_valid & d_first_1;
	wire _T_1211 = ~_T_1005;
	wire _T_1212 = (io_in_d_valid & d_first_1) & ~_T_1005;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [7:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_1005 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [78:0] _GEN_4 = {63'd0, _a_size_lookup_T_5};
	wire [78:0] _d_sizes_clr_T_5 = _GEN_4 << _a_size_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_1211 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1211 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [78:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1211 ? _d_sizes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_1198 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_1222 = inflight >> io_in_d_bits_source;
	wire _T_1224 = _T_1222[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1229 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1230 = (io_in_d_bits_opcode == _GEN_32) | _T_1229;
	wire _T_1234 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1241 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1242 = (io_in_d_bits_opcode == _GEN_48) | _T_1241;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_79 = {4'd0, io_in_d_bits_size};
	wire _T_1246 = _GEN_79 == a_size_lookup;
	wire _T_1256 = (((_T_1209 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_1211;
	wire _T_1258 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set_wo_ready = _GEN_15[4:0];
	wire [4:0] d_clr_wo_ready = _GEN_21[4:0];
	wire _T_1265 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [39:0] a_sizes_set = _GEN_20[39:0];
	wire [39:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [39:0] d_sizes_clr = _GEN_24[39:0];
	wire [39:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [39:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1274 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [39:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [39:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T;
	wire [39:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_75;
	wire [39:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[39:1]};
	wire _T_1300 = (io_in_d_valid & d_first_2) & _T_1005;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_1005 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_1005 ? _d_sizes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_1308 = inflight_1 >> io_in_d_bits_source;
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1318 = _GEN_79 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [39:0] d_sizes_clr_1 = _GEN_69[39:0];
	wire [39:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [39:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	reg [31:0] watchdog_1;
	wire _T_1343 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 40'h0000000000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 40'h0000000000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLAtomicAutomata_1 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [31:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [3:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	reg [1:0] cam_s_0_state;
	reg [2:0] cam_a_0_bits_opcode;
	reg [2:0] cam_a_0_bits_param;
	reg [3:0] cam_a_0_bits_size;
	reg [2:0] cam_a_0_bits_source;
	reg [31:0] cam_a_0_bits_address;
	reg [3:0] cam_a_0_bits_mask;
	reg [31:0] cam_a_0_bits_data;
	reg cam_a_0_bits_corrupt;
	reg [3:0] cam_a_0_lut;
	reg [31:0] cam_d_0_data;
	reg cam_d_0_denied;
	reg cam_d_0_corrupt;
	wire cam_free_0 = cam_s_0_state == 2'h0;
	wire cam_amo_0 = cam_s_0_state == 2'h2;
	wire cam_abusy_0 = (cam_s_0_state == 2'h3) | cam_amo_0;
	wire cam_dmatch_0 = cam_s_0_state != 2'h0;
	wire _a_canLogical_T_1 = auto_in_a_bits_size <= 4'h2;
	wire [31:0] _a_canLogical_T_4 = auto_in_a_bits_address ^ 32'h00002000;
	wire [32:0] _a_canLogical_T_5 = {1'b0, $signed(_a_canLogical_T_4)};
	wire [32:0] _a_canLogical_T_7 = $signed(_a_canLogical_T_5) & 33'sh09a136000;
	wire _a_canLogical_T_8 = $signed(_a_canLogical_T_7) == 33'sh000000000;
	wire [31:0] _a_canLogical_T_9 = auto_in_a_bits_address ^ 32'h00004000;
	wire [32:0] _a_canLogical_T_10 = {1'b0, $signed(_a_canLogical_T_9)};
	wire [32:0] _a_canLogical_T_12 = $signed(_a_canLogical_T_10) & 33'sh09a136000;
	wire _a_canLogical_T_13 = $signed(_a_canLogical_T_12) == 33'sh000000000;
	wire [31:0] _a_canLogical_T_14 = auto_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _a_canLogical_T_15 = {1'b0, $signed(_a_canLogical_T_14)};
	wire [32:0] _a_canLogical_T_17 = $signed(_a_canLogical_T_15) & 33'sh09a136000;
	wire _a_canLogical_T_18 = $signed(_a_canLogical_T_17) == 33'sh000000000;
	wire _a_canLogical_T_20 = (_a_canLogical_T_8 | _a_canLogical_T_13) | _a_canLogical_T_18;
	wire _a_canLogical_T_21 = _a_canLogical_T_1 & _a_canLogical_T_20;
	wire _a_canLogical_T_59 = 4'h2 == auto_in_a_bits_size;
	wire [31:0] _a_canLogical_T_61 = auto_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _a_canLogical_T_62 = {1'b0, $signed(_a_canLogical_T_61)};
	wire [32:0] _a_canLogical_T_64 = $signed(_a_canLogical_T_62) & 33'sh09a134000;
	wire _a_canLogical_T_65 = $signed(_a_canLogical_T_64) == 33'sh000000000;
	wire _a_canLogical_T_66 = _a_canLogical_T_59 & _a_canLogical_T_65;
	wire a_canLogical = _a_canLogical_T_21 | _a_canLogical_T_66;
	wire a_isLogical = auto_in_a_bits_opcode == 3'h3;
	wire a_isArithmetic = auto_in_a_bits_opcode == 3'h2;
	wire _a_isSupported_T = (a_isArithmetic ? a_canLogical : 1'h1);
	wire a_isSupported = (a_isLogical ? a_canLogical : _a_isSupported_T);
	wire [1:0] indexes_0 = {cam_a_0_bits_data[0], cam_d_0_data[0]};
	wire [1:0] indexes_1 = {cam_a_0_bits_data[1], cam_d_0_data[1]};
	wire [1:0] indexes_2 = {cam_a_0_bits_data[2], cam_d_0_data[2]};
	wire [1:0] indexes_3 = {cam_a_0_bits_data[3], cam_d_0_data[3]};
	wire [1:0] indexes_4 = {cam_a_0_bits_data[4], cam_d_0_data[4]};
	wire [1:0] indexes_5 = {cam_a_0_bits_data[5], cam_d_0_data[5]};
	wire [1:0] indexes_6 = {cam_a_0_bits_data[6], cam_d_0_data[6]};
	wire [1:0] indexes_7 = {cam_a_0_bits_data[7], cam_d_0_data[7]};
	wire [1:0] indexes_8 = {cam_a_0_bits_data[8], cam_d_0_data[8]};
	wire [1:0] indexes_9 = {cam_a_0_bits_data[9], cam_d_0_data[9]};
	wire [1:0] indexes_10 = {cam_a_0_bits_data[10], cam_d_0_data[10]};
	wire [1:0] indexes_11 = {cam_a_0_bits_data[11], cam_d_0_data[11]};
	wire [1:0] indexes_12 = {cam_a_0_bits_data[12], cam_d_0_data[12]};
	wire [1:0] indexes_13 = {cam_a_0_bits_data[13], cam_d_0_data[13]};
	wire [1:0] indexes_14 = {cam_a_0_bits_data[14], cam_d_0_data[14]};
	wire [1:0] indexes_15 = {cam_a_0_bits_data[15], cam_d_0_data[15]};
	wire [1:0] indexes_16 = {cam_a_0_bits_data[16], cam_d_0_data[16]};
	wire [1:0] indexes_17 = {cam_a_0_bits_data[17], cam_d_0_data[17]};
	wire [1:0] indexes_18 = {cam_a_0_bits_data[18], cam_d_0_data[18]};
	wire [1:0] indexes_19 = {cam_a_0_bits_data[19], cam_d_0_data[19]};
	wire [1:0] indexes_20 = {cam_a_0_bits_data[20], cam_d_0_data[20]};
	wire [1:0] indexes_21 = {cam_a_0_bits_data[21], cam_d_0_data[21]};
	wire [1:0] indexes_22 = {cam_a_0_bits_data[22], cam_d_0_data[22]};
	wire [1:0] indexes_23 = {cam_a_0_bits_data[23], cam_d_0_data[23]};
	wire [1:0] indexes_24 = {cam_a_0_bits_data[24], cam_d_0_data[24]};
	wire [1:0] indexes_25 = {cam_a_0_bits_data[25], cam_d_0_data[25]};
	wire [1:0] indexes_26 = {cam_a_0_bits_data[26], cam_d_0_data[26]};
	wire [1:0] indexes_27 = {cam_a_0_bits_data[27], cam_d_0_data[27]};
	wire [1:0] indexes_28 = {cam_a_0_bits_data[28], cam_d_0_data[28]};
	wire [1:0] indexes_29 = {cam_a_0_bits_data[29], cam_d_0_data[29]};
	wire [1:0] indexes_30 = {cam_a_0_bits_data[30], cam_d_0_data[30]};
	wire [1:0] indexes_31 = {cam_a_0_bits_data[31], cam_d_0_data[31]};
	wire [3:0] _logic_out_T = cam_a_0_lut >> indexes_0;
	wire [3:0] _logic_out_T_2 = cam_a_0_lut >> indexes_1;
	wire [3:0] _logic_out_T_4 = cam_a_0_lut >> indexes_2;
	wire [3:0] _logic_out_T_6 = cam_a_0_lut >> indexes_3;
	wire [3:0] _logic_out_T_8 = cam_a_0_lut >> indexes_4;
	wire [3:0] _logic_out_T_10 = cam_a_0_lut >> indexes_5;
	wire [3:0] _logic_out_T_12 = cam_a_0_lut >> indexes_6;
	wire [3:0] _logic_out_T_14 = cam_a_0_lut >> indexes_7;
	wire [3:0] _logic_out_T_16 = cam_a_0_lut >> indexes_8;
	wire [3:0] _logic_out_T_18 = cam_a_0_lut >> indexes_9;
	wire [3:0] _logic_out_T_20 = cam_a_0_lut >> indexes_10;
	wire [3:0] _logic_out_T_22 = cam_a_0_lut >> indexes_11;
	wire [3:0] _logic_out_T_24 = cam_a_0_lut >> indexes_12;
	wire [3:0] _logic_out_T_26 = cam_a_0_lut >> indexes_13;
	wire [3:0] _logic_out_T_28 = cam_a_0_lut >> indexes_14;
	wire [3:0] _logic_out_T_30 = cam_a_0_lut >> indexes_15;
	wire [3:0] _logic_out_T_32 = cam_a_0_lut >> indexes_16;
	wire [3:0] _logic_out_T_34 = cam_a_0_lut >> indexes_17;
	wire [3:0] _logic_out_T_36 = cam_a_0_lut >> indexes_18;
	wire [3:0] _logic_out_T_38 = cam_a_0_lut >> indexes_19;
	wire [3:0] _logic_out_T_40 = cam_a_0_lut >> indexes_20;
	wire [3:0] _logic_out_T_42 = cam_a_0_lut >> indexes_21;
	wire [3:0] _logic_out_T_44 = cam_a_0_lut >> indexes_22;
	wire [3:0] _logic_out_T_46 = cam_a_0_lut >> indexes_23;
	wire [3:0] _logic_out_T_48 = cam_a_0_lut >> indexes_24;
	wire [3:0] _logic_out_T_50 = cam_a_0_lut >> indexes_25;
	wire [3:0] _logic_out_T_52 = cam_a_0_lut >> indexes_26;
	wire [3:0] _logic_out_T_54 = cam_a_0_lut >> indexes_27;
	wire [3:0] _logic_out_T_56 = cam_a_0_lut >> indexes_28;
	wire [3:0] _logic_out_T_58 = cam_a_0_lut >> indexes_29;
	wire [3:0] _logic_out_T_60 = cam_a_0_lut >> indexes_30;
	wire [3:0] _logic_out_T_62 = cam_a_0_lut >> indexes_31;
	wire [7:0] logic_out_lo_lo = {_logic_out_T_14[0], _logic_out_T_12[0], _logic_out_T_10[0], _logic_out_T_8[0], _logic_out_T_6[0], _logic_out_T_4[0], _logic_out_T_2[0], _logic_out_T[0]};
	wire [15:0] logic_out_lo = {_logic_out_T_30[0], _logic_out_T_28[0], _logic_out_T_26[0], _logic_out_T_24[0], _logic_out_T_22[0], _logic_out_T_20[0], _logic_out_T_18[0], _logic_out_T_16[0], logic_out_lo_lo};
	wire [7:0] logic_out_hi_lo = {_logic_out_T_46[0], _logic_out_T_44[0], _logic_out_T_42[0], _logic_out_T_40[0], _logic_out_T_38[0], _logic_out_T_36[0], _logic_out_T_34[0], _logic_out_T_32[0]};
	wire [31:0] logic_out = {_logic_out_T_62[0], _logic_out_T_60[0], _logic_out_T_58[0], _logic_out_T_56[0], _logic_out_T_54[0], _logic_out_T_52[0], _logic_out_T_50[0], _logic_out_T_48[0], logic_out_hi_lo, logic_out_lo};
	wire unsigned_ = cam_a_0_bits_param[1];
	wire take_max = cam_a_0_bits_param[0];
	wire adder = cam_a_0_bits_param[2];
	wire [3:0] _signSel_T = ~cam_a_0_bits_mask;
	wire [3:0] _GEN_39 = {1'd0, cam_a_0_bits_mask[3:1]};
	wire [3:0] _signSel_T_2 = _signSel_T | _GEN_39;
	wire [3:0] signSel = ~_signSel_T_2;
	wire [3:0] signbits_a = {cam_a_0_bits_data[31], cam_a_0_bits_data[23], cam_a_0_bits_data[15], cam_a_0_bits_data[7]};
	wire [3:0] signbits_d = {cam_d_0_data[31], cam_d_0_data[23], cam_d_0_data[15], cam_d_0_data[7]};
	wire [3:0] _signbit_a_T = signbits_a & signSel;
	wire [4:0] _signbit_a_T_1 = {_signbit_a_T, 1'h0};
	wire [3:0] signbit_a = _signbit_a_T_1[3:0];
	wire [3:0] _signbit_d_T = signbits_d & signSel;
	wire [4:0] _signbit_d_T_1 = {_signbit_d_T, 1'h0};
	wire [3:0] signbit_d = _signbit_d_T_1[3:0];
	wire [4:0] _signext_a_T = {signbit_a, 1'h0};
	wire [3:0] _signext_a_T_2 = signbit_a | _signext_a_T[3:0];
	wire [5:0] _signext_a_T_3 = {_signext_a_T_2, 2'h0};
	wire [3:0] _signext_a_T_5 = _signext_a_T_2 | _signext_a_T_3[3:0];
	wire [7:0] _signext_a_T_12 = (_signext_a_T_5[0] ? 8'hff : 8'h00);
	wire [7:0] _signext_a_T_14 = (_signext_a_T_5[1] ? 8'hff : 8'h00);
	wire [7:0] _signext_a_T_16 = (_signext_a_T_5[2] ? 8'hff : 8'h00);
	wire [7:0] _signext_a_T_18 = (_signext_a_T_5[3] ? 8'hff : 8'h00);
	wire [31:0] signext_a = {_signext_a_T_18, _signext_a_T_16, _signext_a_T_14, _signext_a_T_12};
	wire [4:0] _signext_d_T = {signbit_d, 1'h0};
	wire [3:0] _signext_d_T_2 = signbit_d | _signext_d_T[3:0];
	wire [5:0] _signext_d_T_3 = {_signext_d_T_2, 2'h0};
	wire [3:0] _signext_d_T_5 = _signext_d_T_2 | _signext_d_T_3[3:0];
	wire [7:0] _signext_d_T_12 = (_signext_d_T_5[0] ? 8'hff : 8'h00);
	wire [7:0] _signext_d_T_14 = (_signext_d_T_5[1] ? 8'hff : 8'h00);
	wire [7:0] _signext_d_T_16 = (_signext_d_T_5[2] ? 8'hff : 8'h00);
	wire [7:0] _signext_d_T_18 = (_signext_d_T_5[3] ? 8'hff : 8'h00);
	wire [31:0] signext_d = {_signext_d_T_18, _signext_d_T_16, _signext_d_T_14, _signext_d_T_12};
	wire [7:0] _wide_mask_T_5 = (cam_a_0_bits_mask[0] ? 8'hff : 8'h00);
	wire [7:0] _wide_mask_T_7 = (cam_a_0_bits_mask[1] ? 8'hff : 8'h00);
	wire [7:0] _wide_mask_T_9 = (cam_a_0_bits_mask[2] ? 8'hff : 8'h00);
	wire [7:0] _wide_mask_T_11 = (cam_a_0_bits_mask[3] ? 8'hff : 8'h00);
	wire [31:0] wide_mask = {_wide_mask_T_11, _wide_mask_T_9, _wide_mask_T_7, _wide_mask_T_5};
	wire [31:0] _a_a_ext_T = cam_a_0_bits_data & wide_mask;
	wire [31:0] a_a_ext = _a_a_ext_T | signext_a;
	wire [31:0] _a_d_ext_T = cam_d_0_data & wide_mask;
	wire [31:0] a_d_ext = _a_d_ext_T | signext_d;
	wire [31:0] _a_d_inv_T = ~a_d_ext;
	wire [31:0] a_d_inv = (adder ? a_d_ext : _a_d_inv_T);
	wire [31:0] adder_out = a_a_ext + a_d_inv;
	wire a_bigger_uneq = unsigned_ == a_a_ext[31];
	wire a_bigger = (a_a_ext[31] == a_d_ext[31] ? ~adder_out[31] : a_bigger_uneq);
	wire pick_a = take_max == a_bigger;
	wire [31:0] _arith_out_T = (pick_a ? cam_a_0_bits_data : cam_d_0_data);
	wire [31:0] arith_out = (adder ? adder_out : _arith_out_T);
	wire [31:0] amo_data = (cam_a_0_bits_opcode[0] ? logic_out : arith_out);
	wire a_allow = ~cam_abusy_0 & (a_isSupported | cam_free_0);
	reg [9:0] beatsLeft;
	wire idle = beatsLeft == 10'h000;
	wire source_i_valid = auto_in_a_valid & a_allow;
	wire [1:0] _readys_T = {source_i_valid, cam_amo_0};
	wire [2:0] _readys_T_1 = {_readys_T, 1'h0};
	wire [1:0] _readys_T_3 = _readys_T | _readys_T_1[1:0];
	wire [2:0] _readys_T_5 = {_readys_T_3, 1'h0};
	wire [1:0] _readys_T_7 = ~_readys_T_5[1:0];
	wire readys_1 = _readys_T_7[1];
	reg state_1;
	wire allowed_1 = (idle ? readys_1 : state_1);
	wire out_1_ready = auto_out_a_ready & allowed_1;
	wire _T = ~a_isSupported;
	wire [2:0] source_i_bits_opcode = (~a_isSupported ? 3'h4 : auto_in_a_bits_opcode);
	wire [2:0] source_i_bits_param = (~a_isSupported ? 3'h0 : auto_in_a_bits_param);
	wire source_c_bits_a_corrupt = cam_a_0_bits_corrupt | cam_d_0_corrupt;
	wire source_c_bits_a_mask_sizeOH_shiftAmount = cam_a_0_bits_size[0];
	wire [1:0] _source_c_bits_a_mask_sizeOH_T_1 = 2'h1 << source_c_bits_a_mask_sizeOH_shiftAmount;
	wire [1:0] source_c_bits_a_mask_sizeOH = _source_c_bits_a_mask_sizeOH_T_1 | 2'h1;
	wire _source_c_bits_a_mask_T = cam_a_0_bits_size >= 4'h2;
	wire source_c_bits_a_mask_size = source_c_bits_a_mask_sizeOH[1];
	wire source_c_bits_a_mask_bit = cam_a_0_bits_address[1];
	wire source_c_bits_a_mask_nbit = ~source_c_bits_a_mask_bit;
	wire source_c_bits_a_mask_acc = _source_c_bits_a_mask_T | (source_c_bits_a_mask_size & source_c_bits_a_mask_nbit);
	wire source_c_bits_a_mask_acc_1 = _source_c_bits_a_mask_T | (source_c_bits_a_mask_size & source_c_bits_a_mask_bit);
	wire source_c_bits_a_mask_size_1 = source_c_bits_a_mask_sizeOH[0];
	wire source_c_bits_a_mask_bit_1 = cam_a_0_bits_address[0];
	wire source_c_bits_a_mask_nbit_1 = ~source_c_bits_a_mask_bit_1;
	wire source_c_bits_a_mask_eq_2 = source_c_bits_a_mask_nbit & source_c_bits_a_mask_nbit_1;
	wire source_c_bits_a_mask_acc_2 = source_c_bits_a_mask_acc | (source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_2);
	wire source_c_bits_a_mask_eq_3 = source_c_bits_a_mask_nbit & source_c_bits_a_mask_bit_1;
	wire source_c_bits_a_mask_acc_3 = source_c_bits_a_mask_acc | (source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_3);
	wire source_c_bits_a_mask_eq_4 = source_c_bits_a_mask_bit & source_c_bits_a_mask_nbit_1;
	wire source_c_bits_a_mask_acc_4 = source_c_bits_a_mask_acc_1 | (source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_4);
	wire source_c_bits_a_mask_eq_5 = source_c_bits_a_mask_bit & source_c_bits_a_mask_bit_1;
	wire source_c_bits_a_mask_acc_5 = source_c_bits_a_mask_acc_1 | (source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_5);
	wire [3:0] source_c_bits_a_mask = {source_c_bits_a_mask_acc_5, source_c_bits_a_mask_acc_4, source_c_bits_a_mask_acc_3, source_c_bits_a_mask_acc_2};
	wire [26:0] _decode_T_1 = 27'h0000fff << auto_in_a_bits_size;
	wire [11:0] _decode_T_3 = ~_decode_T_1[11:0];
	wire [9:0] decode = _decode_T_3[11:2];
	wire opdata = ~auto_in_a_bits_opcode[2];
	wire latch = idle & auto_out_a_ready;
	wire readys_0 = _readys_T_7[0];
	wire earlyWinner_0 = readys_0 & cam_amo_0;
	wire earlyWinner_1 = readys_1 & source_i_valid;
	wire _prefixOR_T = earlyWinner_0 | earlyWinner_1;
	wire _T_10 = ~reset;
	wire _T_12 = cam_amo_0 | source_i_valid;
	wire _T_13 = ~(cam_amo_0 | source_i_valid);
	reg state_0;
	wire muxStateEarly_0 = (idle ? earlyWinner_0 : state_0);
	wire muxStateEarly_1 = (idle ? earlyWinner_1 : state_1);
	wire _sink_ACancel_earlyValid_T_3 = (state_0 & cam_amo_0) | (state_1 & source_i_valid);
	wire sink_ACancel_earlyValid = (idle ? _T_12 : _sink_ACancel_earlyValid_T_3);
	wire _beatsLeft_T_2 = auto_out_a_ready & sink_ACancel_earlyValid;
	wire [9:0] _GEN_40 = {9'd0, _beatsLeft_T_2};
	wire [9:0] _beatsLeft_T_4 = beatsLeft - _GEN_40;
	wire allowed_0 = (idle ? readys_0 : state_0);
	wire out_ready = auto_out_a_ready & allowed_0;
	wire [31:0] _T_29 = (muxStateEarly_0 ? amo_data : 32'h00000000);
	wire [31:0] _T_30 = (muxStateEarly_1 ? auto_in_a_bits_data : 32'h00000000);
	wire [3:0] _T_32 = (muxStateEarly_0 ? source_c_bits_a_mask : 4'h0);
	wire [3:0] _T_33 = (muxStateEarly_1 ? auto_in_a_bits_mask : 4'h0);
	wire [31:0] _T_35 = (muxStateEarly_0 ? cam_a_0_bits_address : 32'h00000000);
	wire [31:0] _T_36 = (muxStateEarly_1 ? auto_in_a_bits_address : 32'h00000000);
	wire [2:0] _T_38 = (muxStateEarly_0 ? cam_a_0_bits_source : 3'h0);
	wire [2:0] _T_39 = (muxStateEarly_1 ? auto_in_a_bits_source : 3'h0);
	wire [3:0] _T_41 = (muxStateEarly_0 ? cam_a_0_bits_size : 4'h0);
	wire [3:0] _T_42 = (muxStateEarly_1 ? auto_in_a_bits_size : 4'h0);
	wire _T_50 = out_1_ready & source_i_valid;
	wire [2:0] _GEN_41 = {1'd0, auto_in_a_bits_param[1:0]};
	wire [3:0] _cam_a_0_lut_T_2 = (3'h1 == _GEN_41 ? 4'he : 4'h8);
	wire [1:0] _GEN_12 = (cam_free_0 ? 2'h3 : cam_s_0_state);
	wire [1:0] _GEN_23 = (_T_50 & _T ? _GEN_12 : cam_s_0_state);
	wire _T_53 = out_ready & cam_amo_0;
	wire [1:0] _GEN_24 = (cam_amo_0 ? 2'h1 : _GEN_23);
	wire [1:0] _GEN_25 = (_T_53 ? _GEN_24 : _GEN_23);
	reg [9:0] d_first_counter;
	wire d_first = d_first_counter == 10'h000;
	wire d_ackd = auto_out_d_bits_opcode == 3'h1;
	wire d_cam_sel_raw_0 = cam_a_0_bits_source == auto_out_d_bits_source;
	wire d_cam_sel_match_0 = d_cam_sel_raw_0 & cam_dmatch_0;
	wire d_drop = (d_first & d_ackd) & d_cam_sel_match_0;
	wire bundleOut_0_d_ready = auto_in_d_ready | d_drop;
	wire _d_first_T = bundleOut_0_d_ready & auto_out_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << auto_out_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = auto_out_d_bits_opcode[0];
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_ack = auto_out_d_bits_opcode == 3'h0;
	wire d_replace = (d_first & d_ack) & d_cam_sel_match_0;
	TLMonitor_20 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	assign auto_in_a_ready = out_1_ready & a_allow;
	assign auto_in_d_valid = auto_out_d_valid & ~d_drop;
	assign auto_in_d_bits_opcode = (d_replace ? 3'h1 : auto_out_d_bits_opcode);
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = (d_replace ? cam_d_0_denied | auto_out_d_bits_denied : auto_out_d_bits_denied);
	assign auto_in_d_bits_data = (d_replace ? cam_d_0_data : auto_out_d_bits_data);
	assign auto_in_d_bits_corrupt = (d_replace ? cam_d_0_corrupt | auto_out_d_bits_denied : auto_out_d_bits_corrupt);
	assign auto_out_a_valid = (idle ? _T_12 : _sink_ACancel_earlyValid_T_3);
	assign auto_out_a_bits_opcode = (muxStateEarly_1 ? source_i_bits_opcode : 3'h0);
	assign auto_out_a_bits_param = (muxStateEarly_1 ? source_i_bits_param : 3'h0);
	assign auto_out_a_bits_size = _T_41 | _T_42;
	assign auto_out_a_bits_source = _T_38 | _T_39;
	assign auto_out_a_bits_address = _T_35 | _T_36;
	assign auto_out_a_bits_mask = _T_32 | _T_33;
	assign auto_out_a_bits_data = _T_29 | _T_30;
	assign auto_out_a_bits_corrupt = (muxStateEarly_0 & source_c_bits_a_corrupt) | (muxStateEarly_1 & auto_in_a_bits_corrupt);
	assign auto_out_d_ready = auto_in_d_ready | d_drop;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = out_1_ready & a_allow;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid & ~d_drop;
	assign monitor_io_in_d_bits_opcode = (d_replace ? 3'h1 : auto_out_d_bits_opcode);
	assign monitor_io_in_d_bits_param = auto_out_d_bits_param;
	assign monitor_io_in_d_bits_size = auto_out_d_bits_size;
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source;
	assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink;
	assign monitor_io_in_d_bits_denied = (d_replace ? cam_d_0_denied | auto_out_d_bits_denied : auto_out_d_bits_denied);
	assign monitor_io_in_d_bits_corrupt = (d_replace ? cam_d_0_corrupt | auto_out_d_bits_denied : auto_out_d_bits_corrupt);
	always @(posedge clock) begin
		if (reset)
			cam_s_0_state <= 2'h0;
		else if (_d_first_T & d_first) begin
			if (d_cam_sel_match_0) begin
				if (d_ackd)
					cam_s_0_state <= 2'h2;
				else
					cam_s_0_state <= 2'h0;
			end
			else
				cam_s_0_state <= _GEN_25;
		end
		else
			cam_s_0_state <= _GEN_25;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_opcode <= auto_in_a_bits_opcode;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_param <= auto_in_a_bits_param;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_size <= auto_in_a_bits_size;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_source <= auto_in_a_bits_source;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_address <= auto_in_a_bits_address;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_mask <= auto_in_a_bits_mask;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_data <= auto_in_a_bits_data;
		if (_T_50 & _T)
			if (cam_free_0)
				cam_a_0_bits_corrupt <= auto_in_a_bits_corrupt;
		if (_T_50 & _T)
			if (cam_free_0)
				if (3'h3 == _GEN_41)
					cam_a_0_lut <= 4'hc;
				else if (3'h0 == _GEN_41)
					cam_a_0_lut <= 4'h6;
				else
					cam_a_0_lut <= _cam_a_0_lut_T_2;
		if (_d_first_T & d_first)
			if (d_cam_sel_match_0 & d_ackd)
				cam_d_0_data <= auto_out_d_bits_data;
		if (_d_first_T & d_first)
			if (d_cam_sel_match_0 & d_ackd)
				cam_d_0_denied <= auto_out_d_bits_denied;
		if (_d_first_T & d_first)
			if (d_cam_sel_match_0 & d_ackd)
				cam_d_0_corrupt <= auto_out_d_bits_corrupt;
		if (reset)
			beatsLeft <= 10'h000;
		else if (latch) begin
			if (earlyWinner_1) begin
				if (opdata)
					beatsLeft <= decode;
				else
					beatsLeft <= 10'h000;
			end
			else
				beatsLeft <= 10'h000;
		end
		else
			beatsLeft <= _beatsLeft_T_4;
		if (reset)
			state_1 <= 1'h0;
		else if (idle)
			state_1 <= earlyWinner_1;
		if (reset)
			state_0 <= 1'h0;
		else if (idle)
			state_0 <= earlyWinner_0;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
	end
endmodule
module TLMonitor_21 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [13:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [3:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [13:0] _GEN_71 = {2'd0, is_aligned_mask};
	wire [13:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 14'h0000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire _T_44 = io_in_a_bits_size <= 4'hc;
	wire _T_53 = _T_44 & source_ok;
	wire [13:0] _T_56 = io_in_a_bits_address ^ 14'h3000;
	wire [14:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [14:0] _T_59 = $signed(_T_57) & -15'sh1000;
	wire _T_60 = $signed(_T_59) == 15'sh0000;
	wire _T_76 = _T_44 & _T_60;
	wire _T_92 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_96 = ~io_in_a_bits_mask;
	wire _T_97 = _T_96 == 4'h0;
	wire _T_101 = ~io_in_a_bits_corrupt;
	wire _T_105 = io_in_a_bits_opcode == 3'h7;
	wire _T_159 = io_in_a_bits_param != 3'h0;
	wire _T_172 = io_in_a_bits_opcode == 3'h4;
	wire _T_208 = io_in_a_bits_param == 3'h0;
	wire _T_212 = io_in_a_bits_mask == mask;
	wire _T_220 = io_in_a_bits_opcode == 3'h0;
	wire _T_244 = _T_53 & _T_76;
	wire _T_262 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_300 = ~mask;
	wire [3:0] _T_301 = io_in_a_bits_mask & _T_300;
	wire _T_302 = _T_301 == 4'h0;
	wire _T_306 = io_in_a_bits_opcode == 3'h2;
	wire _T_320 = io_in_a_bits_size <= 4'h2;
	wire _T_328 = _T_320 & _T_60;
	wire _T_330 = _T_53 & _T_328;
	wire _T_340 = io_in_a_bits_param <= 3'h4;
	wire _T_348 = io_in_a_bits_opcode == 3'h3;
	wire _T_382 = io_in_a_bits_param <= 3'h3;
	wire _T_390 = io_in_a_bits_opcode == 3'h5;
	wire _T_424 = io_in_a_bits_param <= 3'h1;
	wire _T_436 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_440 = io_in_d_bits_opcode == 3'h6;
	wire _T_444 = io_in_d_bits_size >= 4'h2;
	wire _T_452 = ~io_in_d_bits_corrupt;
	wire _T_460 = io_in_d_bits_opcode == 3'h4;
	wire _T_488 = io_in_d_bits_opcode == 3'h5;
	wire _T_517 = io_in_d_bits_opcode == 3'h0;
	wire _T_534 = io_in_d_bits_opcode == 3'h1;
	wire _T_552 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg [2:0] source;
	reg [13:0] address;
	wire _T_582 = io_in_a_valid & ~a_first;
	wire _T_583 = io_in_a_bits_opcode == opcode;
	wire _T_587 = io_in_a_bits_param == param;
	wire _T_591 = io_in_a_bits_size == size;
	wire _T_595 = io_in_a_bits_source == source;
	wire _T_599 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [3:0] size_1;
	reg [2:0] source_1;
	wire _T_606 = io_in_d_valid & ~d_first;
	wire _T_607 = io_in_d_bits_opcode == opcode_1;
	wire _T_615 = io_in_d_bits_size == size_1;
	wire _T_619 = io_in_d_bits_source == source_1;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [39:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [5:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0};
	wire [39:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T;
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [39:0] _GEN_75 = {24'd0, _a_size_lookup_T_5};
	wire [39:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_75;
	wire [39:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[39:1]};
	wire _T_633 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire [7:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire _T_636 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [4:0] _GEN_77 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_77};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [5:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [67:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [67:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire [4:0] _T_638 = inflight >> io_in_a_bits_source;
	wire _T_640 = ~_T_638[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [67:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 68'h00000000000000000);
	wire _T_644 = io_in_d_valid & d_first_1;
	wire _T_646 = ~_T_440;
	wire _T_647 = (io_in_d_valid & d_first_1) & ~_T_440;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [7:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_440 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [78:0] _GEN_4 = {63'd0, _a_size_lookup_T_5};
	wire [78:0] _d_sizes_clr_T_5 = _GEN_4 << _a_size_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_646 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_646 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [78:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_646 ? _d_sizes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_633 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_657 = inflight >> io_in_d_bits_source;
	wire _T_659 = _T_657[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_664 = io_in_d_bits_opcode == _GEN_40;
	wire _T_665 = (io_in_d_bits_opcode == _GEN_32) | _T_664;
	wire _T_669 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_676 = io_in_d_bits_opcode == _GEN_56;
	wire _T_677 = (io_in_d_bits_opcode == _GEN_48) | _T_676;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_79 = {4'd0, io_in_d_bits_size};
	wire _T_681 = _GEN_79 == a_size_lookup;
	wire _T_691 = (((_T_644 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_646;
	wire _T_693 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set_wo_ready = _GEN_15[4:0];
	wire [4:0] d_clr_wo_ready = _GEN_21[4:0];
	wire _T_700 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [39:0] a_sizes_set = _GEN_20[39:0];
	wire [39:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [39:0] d_sizes_clr = _GEN_24[39:0];
	wire [39:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [39:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_709 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [39:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [39:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T;
	wire [39:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_75;
	wire [39:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[39:1]};
	wire _T_735 = (io_in_d_valid & d_first_2) & _T_440;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_440 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_440 ? _d_sizes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_743 = inflight_1 >> io_in_d_bits_source;
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_753 = _GEN_79 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [39:0] d_sizes_clr_1 = _GEN_69[39:0];
	wire [39:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [39:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	reg [31:0] watchdog_1;
	wire _T_778 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 40'h0000000000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 40'h0000000000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Queue_10 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_size,
	io_enq_bits_source,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_size,
	io_deq_bits_source
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [3:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [3:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	reg [2:0] ram_opcode [0:0];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [3:0] ram_size [0:0];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [3:0] ram_size_io_deq_bits_MPORT_data;
	wire [3:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg [2:0] ram_source [0:0];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire [2:0] ram_source_io_deq_bits_MPORT_data;
	wire [2:0] ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg maybe_full;
	wire empty = ~maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = 1'h0;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = 1'h0;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = 1'h0;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = 1'h0;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = 1'h0;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~maybe_full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module TLError (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [13:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [3:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [13:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [3:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_corrupt;
	wire a_clock;
	wire a_reset;
	wire a_io_enq_ready;
	wire a_io_enq_valid;
	wire [2:0] a_io_enq_bits_opcode;
	wire [3:0] a_io_enq_bits_size;
	wire [2:0] a_io_enq_bits_source;
	wire a_io_deq_ready;
	wire a_io_deq_valid;
	wire [2:0] a_io_deq_bits_opcode;
	wire [3:0] a_io_deq_bits_size;
	wire [2:0] a_io_deq_bits_source;
	wire _a_last_T = a_io_deq_ready & a_io_deq_valid;
	wire [26:0] _a_last_beats1_decode_T_1 = 27'h0000fff << a_io_deq_bits_size;
	wire [11:0] _a_last_beats1_decode_T_3 = ~_a_last_beats1_decode_T_1[11:0];
	wire [9:0] a_last_beats1_decode = _a_last_beats1_decode_T_3[11:2];
	wire a_last_beats1_opdata = ~a_io_deq_bits_opcode[2];
	wire [9:0] a_last_beats1 = (a_last_beats1_opdata ? a_last_beats1_decode : 10'h000);
	reg [9:0] a_last_counter;
	wire [9:0] a_last_counter1 = a_last_counter - 10'h001;
	wire a_last_first = a_last_counter == 10'h000;
	wire a_last = (a_last_counter == 10'h001) | (a_last_beats1 == 10'h000);
	wire da_valid = a_io_deq_valid & a_last;
	wire _T = auto_in_d_ready & da_valid;
	wire [3:0] da_bits_size = a_io_deq_bits_size;
	wire [26:0] _beats1_decode_T_1 = 27'h0000fff << da_bits_size;
	wire [11:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[11:0];
	wire [9:0] beats1_decode = _beats1_decode_T_3[11:2];
	wire [2:0] _GEN_4 = (3'h2 == a_io_deq_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_5 = (3'h3 == a_io_deq_bits_opcode ? 3'h1 : _GEN_4);
	wire [2:0] _GEN_6 = (3'h4 == a_io_deq_bits_opcode ? 3'h1 : _GEN_5);
	wire [2:0] _GEN_7 = (3'h5 == a_io_deq_bits_opcode ? 3'h2 : _GEN_6);
	wire [2:0] _GEN_8 = (3'h6 == a_io_deq_bits_opcode ? 3'h4 : _GEN_7);
	wire [2:0] da_bits_opcode = (3'h7 == a_io_deq_bits_opcode ? 3'h4 : _GEN_8);
	wire beats1_opdata = da_bits_opcode[0];
	wire [9:0] beats1 = (beats1_opdata ? beats1_decode : 10'h000);
	reg [9:0] counter;
	wire [9:0] counter1 = counter - 10'h001;
	wire da_first = counter == 10'h000;
	wire da_last = (counter == 10'h001) | (beats1 == 10'h000);
	TLMonitor_21 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Queue_10 a(
		.clock(a_clock),
		.reset(a_reset),
		.io_enq_ready(a_io_enq_ready),
		.io_enq_valid(a_io_enq_valid),
		.io_enq_bits_opcode(a_io_enq_bits_opcode),
		.io_enq_bits_size(a_io_enq_bits_size),
		.io_enq_bits_source(a_io_enq_bits_source),
		.io_deq_ready(a_io_deq_ready),
		.io_deq_valid(a_io_deq_valid),
		.io_deq_bits_opcode(a_io_deq_bits_opcode),
		.io_deq_bits_size(a_io_deq_bits_size),
		.io_deq_bits_source(a_io_deq_bits_source)
	);
	assign auto_in_a_ready = a_io_enq_ready;
	assign auto_in_d_valid = a_io_deq_valid & a_last;
	assign auto_in_d_bits_opcode = (3'h7 == a_io_deq_bits_opcode ? 3'h4 : _GEN_8);
	assign auto_in_d_bits_size = a_io_deq_bits_size;
	assign auto_in_d_bits_source = a_io_deq_bits_source;
	assign auto_in_d_bits_corrupt = da_bits_opcode[0];
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = a_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = a_io_deq_valid & a_last;
	assign monitor_io_in_d_bits_opcode = (3'h7 == a_io_deq_bits_opcode ? 3'h4 : _GEN_8);
	assign monitor_io_in_d_bits_size = a_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = a_io_deq_bits_source;
	assign monitor_io_in_d_bits_corrupt = da_bits_opcode[0];
	assign a_clock = clock;
	assign a_reset = reset;
	assign a_io_enq_valid = auto_in_a_valid;
	assign a_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign a_io_enq_bits_size = auto_in_a_bits_size;
	assign a_io_enq_bits_source = auto_in_a_bits_source;
	assign a_io_deq_ready = (auto_in_d_ready & da_last) | ~a_last;
	always @(posedge clock) begin
		if (reset)
			a_last_counter <= 10'h000;
		else if (_a_last_T)
			if (a_last_first) begin
				if (a_last_beats1_opdata)
					a_last_counter <= a_last_beats1_decode;
				else
					a_last_counter <= 10'h000;
			end
			else
				a_last_counter <= a_last_counter1;
		if (reset)
			counter <= 10'h000;
		else if (_T)
			if (da_first) begin
				if (beats1_opdata)
					counter <= beats1_decode;
				else
					counter <= 10'h000;
			end
			else
				counter <= counter1;
	end
endmodule
module TLMonitor_22 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [13:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [13:0] _GEN_71 = {2'd0, is_aligned_mask};
	wire [13:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 14'h0000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire _T_44 = io_in_a_bits_size <= 4'hc;
	wire _T_53 = _T_44 & source_ok;
	wire [13:0] _T_56 = io_in_a_bits_address ^ 14'h3000;
	wire [14:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [14:0] _T_59 = $signed(_T_57) & -15'sh1000;
	wire _T_60 = $signed(_T_59) == 15'sh0000;
	wire _T_76 = _T_44 & _T_60;
	wire _T_92 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_96 = ~io_in_a_bits_mask;
	wire _T_97 = _T_96 == 4'h0;
	wire _T_101 = ~io_in_a_bits_corrupt;
	wire _T_105 = io_in_a_bits_opcode == 3'h7;
	wire _T_159 = io_in_a_bits_param != 3'h0;
	wire _T_172 = io_in_a_bits_opcode == 3'h4;
	wire _T_208 = io_in_a_bits_param == 3'h0;
	wire _T_212 = io_in_a_bits_mask == mask;
	wire _T_220 = io_in_a_bits_opcode == 3'h0;
	wire _T_244 = _T_53 & _T_76;
	wire _T_262 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_300 = ~mask;
	wire [3:0] _T_301 = io_in_a_bits_mask & _T_300;
	wire _T_302 = _T_301 == 4'h0;
	wire _T_306 = io_in_a_bits_opcode == 3'h2;
	wire _T_320 = io_in_a_bits_size <= 4'h2;
	wire _T_328 = _T_320 & _T_60;
	wire _T_330 = _T_53 & _T_328;
	wire _T_340 = io_in_a_bits_param <= 3'h4;
	wire _T_348 = io_in_a_bits_opcode == 3'h3;
	wire _T_382 = io_in_a_bits_param <= 3'h3;
	wire _T_390 = io_in_a_bits_opcode == 3'h5;
	wire _T_424 = io_in_a_bits_param <= 3'h1;
	wire _T_436 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_440 = io_in_d_bits_opcode == 3'h6;
	wire _T_444 = io_in_d_bits_size >= 4'h2;
	wire _T_448 = io_in_d_bits_param == 2'h0;
	wire _T_452 = ~io_in_d_bits_corrupt;
	wire _T_456 = ~io_in_d_bits_denied;
	wire _T_460 = io_in_d_bits_opcode == 3'h4;
	wire _T_471 = io_in_d_bits_param <= 2'h2;
	wire _T_475 = io_in_d_bits_param != 2'h2;
	wire _T_488 = io_in_d_bits_opcode == 3'h5;
	wire _T_508 = _T_456 | io_in_d_bits_corrupt;
	wire _T_517 = io_in_d_bits_opcode == 3'h0;
	wire _T_534 = io_in_d_bits_opcode == 3'h1;
	wire _T_552 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg [2:0] source;
	reg [13:0] address;
	wire _T_582 = io_in_a_valid & ~a_first;
	wire _T_583 = io_in_a_bits_opcode == opcode;
	wire _T_587 = io_in_a_bits_param == param;
	wire _T_591 = io_in_a_bits_size == size;
	wire _T_595 = io_in_a_bits_source == source;
	wire _T_599 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_606 = io_in_d_valid & ~d_first;
	wire _T_607 = io_in_d_bits_opcode == opcode_1;
	wire _T_611 = io_in_d_bits_param == param_1;
	wire _T_615 = io_in_d_bits_size == size_1;
	wire _T_619 = io_in_d_bits_source == source_1;
	wire _T_623 = io_in_d_bits_sink == sink;
	wire _T_627 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [39:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [5:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0};
	wire [39:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T;
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [39:0] _GEN_75 = {24'd0, _a_size_lookup_T_5};
	wire [39:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_75;
	wire [39:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[39:1]};
	wire _T_633 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire [7:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire _T_636 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [4:0] _GEN_77 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_77};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [5:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [67:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [67:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire [4:0] _T_638 = inflight >> io_in_a_bits_source;
	wire _T_640 = ~_T_638[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [67:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 68'h00000000000000000);
	wire _T_644 = io_in_d_valid & d_first_1;
	wire _T_646 = ~_T_440;
	wire _T_647 = (io_in_d_valid & d_first_1) & ~_T_440;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [7:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_440 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [78:0] _GEN_4 = {63'd0, _a_size_lookup_T_5};
	wire [78:0] _d_sizes_clr_T_5 = _GEN_4 << _a_size_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_646 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_646 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [78:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_646 ? _d_sizes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_633 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_657 = inflight >> io_in_d_bits_source;
	wire _T_659 = _T_657[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_664 = io_in_d_bits_opcode == _GEN_40;
	wire _T_665 = (io_in_d_bits_opcode == _GEN_32) | _T_664;
	wire _T_669 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_676 = io_in_d_bits_opcode == _GEN_56;
	wire _T_677 = (io_in_d_bits_opcode == _GEN_48) | _T_676;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_79 = {4'd0, io_in_d_bits_size};
	wire _T_681 = _GEN_79 == a_size_lookup;
	wire _T_691 = (((_T_644 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_646;
	wire _T_693 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set_wo_ready = _GEN_15[4:0];
	wire [4:0] d_clr_wo_ready = _GEN_21[4:0];
	wire _T_700 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [39:0] a_sizes_set = _GEN_20[39:0];
	wire [39:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [39:0] d_sizes_clr = _GEN_24[39:0];
	wire [39:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [39:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_709 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [39:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [39:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T;
	wire [39:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_75;
	wire [39:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[39:1]};
	wire _T_735 = (io_in_d_valid & d_first_2) & _T_440;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_440 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_440 ? _d_sizes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_743 = inflight_1 >> io_in_d_bits_source;
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_753 = _GEN_79 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [39:0] d_sizes_clr_1 = _GEN_69[39:0];
	wire [39:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [39:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	reg [31:0] watchdog_1;
	wire _T_778 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 40'h0000000000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 40'h0000000000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Queue_11 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [3:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [13:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [3:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [13:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire io_deq_bits_corrupt;
	reg [2:0] ram_opcode [0:1];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [2:0] ram_param [0:1];
	wire ram_param_io_deq_bits_MPORT_en;
	wire ram_param_io_deq_bits_MPORT_addr;
	wire [2:0] ram_param_io_deq_bits_MPORT_data;
	wire [2:0] ram_param_MPORT_data;
	wire ram_param_MPORT_addr;
	wire ram_param_MPORT_mask;
	wire ram_param_MPORT_en;
	reg [3:0] ram_size [0:1];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [3:0] ram_size_io_deq_bits_MPORT_data;
	wire [3:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg [2:0] ram_source [0:1];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire [2:0] ram_source_io_deq_bits_MPORT_data;
	wire [2:0] ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg [13:0] ram_address [0:1];
	wire ram_address_io_deq_bits_MPORT_en;
	wire ram_address_io_deq_bits_MPORT_addr;
	wire [13:0] ram_address_io_deq_bits_MPORT_data;
	wire [13:0] ram_address_MPORT_data;
	wire ram_address_MPORT_addr;
	wire ram_address_MPORT_mask;
	wire ram_address_MPORT_en;
	reg [3:0] ram_mask [0:1];
	wire ram_mask_io_deq_bits_MPORT_en;
	wire ram_mask_io_deq_bits_MPORT_addr;
	wire [3:0] ram_mask_io_deq_bits_MPORT_data;
	wire [3:0] ram_mask_MPORT_data;
	wire ram_mask_MPORT_addr;
	wire ram_mask_MPORT_mask;
	wire ram_mask_MPORT_en;
	reg ram_corrupt [0:1];
	wire ram_corrupt_io_deq_bits_MPORT_en;
	wire ram_corrupt_io_deq_bits_MPORT_addr;
	wire ram_corrupt_io_deq_bits_MPORT_data;
	wire ram_corrupt_MPORT_data;
	wire ram_corrupt_MPORT_addr;
	wire ram_corrupt_MPORT_mask;
	wire ram_corrupt_MPORT_en;
	reg value;
	reg value_1;
	reg maybe_full;
	wire ptr_match = value == value_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = value;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_param_io_deq_bits_MPORT_en = 1'h1;
	assign ram_param_io_deq_bits_MPORT_addr = value_1;
	assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr];
	assign ram_param_MPORT_data = io_enq_bits_param;
	assign ram_param_MPORT_addr = value;
	assign ram_param_MPORT_mask = 1'h1;
	assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = value_1;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = value;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = value_1;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = value;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_address_io_deq_bits_MPORT_en = 1'h1;
	assign ram_address_io_deq_bits_MPORT_addr = value_1;
	assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr];
	assign ram_address_MPORT_data = io_enq_bits_address;
	assign ram_address_MPORT_addr = value;
	assign ram_address_MPORT_mask = 1'h1;
	assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
	assign ram_mask_io_deq_bits_MPORT_addr = value_1;
	assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr];
	assign ram_mask_MPORT_data = io_enq_bits_mask;
	assign ram_mask_MPORT_addr = value;
	assign ram_mask_MPORT_mask = 1'h1;
	assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
	assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
	assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr];
	assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
	assign ram_corrupt_MPORT_addr = value;
	assign ram_corrupt_MPORT_mask = 1'h1;
	assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data;
	assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data;
	assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_param_MPORT_en & ram_param_MPORT_mask)
			ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (ram_address_MPORT_en & ram_address_MPORT_mask)
			ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data;
		if (ram_mask_MPORT_en & ram_mask_MPORT_mask)
			ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data;
		if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask)
			ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data;
		if (reset)
			value <= 1'h0;
		else if (do_enq)
			value <= value + 1'h1;
		if (reset)
			value_1 <= 1'h0;
		else if (do_deq)
			value_1 <= value_1 + 1'h1;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module TLBuffer_7 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [13:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [13:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [3:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [13:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [3:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire bundleOut_0_a_q_clock;
	wire bundleOut_0_a_q_reset;
	wire bundleOut_0_a_q_io_enq_ready;
	wire bundleOut_0_a_q_io_enq_valid;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_param;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_size;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_source;
	wire [13:0] bundleOut_0_a_q_io_enq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_mask;
	wire bundleOut_0_a_q_io_enq_bits_corrupt;
	wire bundleOut_0_a_q_io_deq_ready;
	wire bundleOut_0_a_q_io_deq_valid;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_param;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_size;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_source;
	wire [13:0] bundleOut_0_a_q_io_deq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_mask;
	wire bundleOut_0_a_q_io_deq_bits_corrupt;
	wire bundleIn_0_d_q_clock;
	wire bundleIn_0_d_q_reset;
	wire bundleIn_0_d_q_io_enq_ready;
	wire bundleIn_0_d_q_io_enq_valid;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_enq_bits_param;
	wire [3:0] bundleIn_0_d_q_io_enq_bits_size;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_source;
	wire bundleIn_0_d_q_io_enq_bits_sink;
	wire bundleIn_0_d_q_io_enq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_enq_bits_data;
	wire bundleIn_0_d_q_io_enq_bits_corrupt;
	wire bundleIn_0_d_q_io_deq_ready;
	wire bundleIn_0_d_q_io_deq_valid;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_param;
	wire [3:0] bundleIn_0_d_q_io_deq_bits_size;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_source;
	wire bundleIn_0_d_q_io_deq_bits_sink;
	wire bundleIn_0_d_q_io_deq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_deq_bits_data;
	wire bundleIn_0_d_q_io_deq_bits_corrupt;
	TLMonitor_22 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Queue_11 bundleOut_0_a_q(
		.clock(bundleOut_0_a_q_clock),
		.reset(bundleOut_0_a_q_reset),
		.io_enq_ready(bundleOut_0_a_q_io_enq_ready),
		.io_enq_valid(bundleOut_0_a_q_io_enq_valid),
		.io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
		.io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
		.io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
		.io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
		.io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
		.io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleOut_0_a_q_io_deq_ready),
		.io_deq_valid(bundleOut_0_a_q_io_deq_valid),
		.io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
		.io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
		.io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
		.io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
		.io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
		.io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
	);
	Queue_9 bundleIn_0_d_q(
		.clock(bundleIn_0_d_q_clock),
		.reset(bundleIn_0_d_q_reset),
		.io_enq_ready(bundleIn_0_d_q_io_enq_ready),
		.io_enq_valid(bundleIn_0_d_q_io_enq_valid),
		.io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
		.io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
		.io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
		.io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
		.io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
		.io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleIn_0_d_q_io_deq_ready),
		.io_deq_valid(bundleIn_0_d_q_io_deq_valid),
		.io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
		.io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
		.io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
		.io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
		.io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
		.io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data;
	assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid;
	assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode;
	assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param;
	assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size;
	assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source;
	assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address;
	assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask;
	assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt;
	assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign bundleOut_0_a_q_clock = clock;
	assign bundleOut_0_a_q_reset = reset;
	assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid;
	assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param;
	assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size;
	assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source;
	assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address;
	assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask;
	assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready;
	assign bundleIn_0_d_q_clock = clock;
	assign bundleIn_0_d_q_reset = reset;
	assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid;
	assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign bundleIn_0_d_q_io_enq_bits_param = 2'h0;
	assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size;
	assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source;
	assign bundleIn_0_d_q_io_enq_bits_sink = 1'h0;
	assign bundleIn_0_d_q_io_enq_bits_denied = 1'h1;
	assign bundleIn_0_d_q_io_enq_bits_data = 32'h00000000;
	assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt;
	assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready;
endmodule
module ErrorDeviceWrapper (
	clock,
	reset,
	auto_buffer_in_a_ready,
	auto_buffer_in_a_valid,
	auto_buffer_in_a_bits_opcode,
	auto_buffer_in_a_bits_param,
	auto_buffer_in_a_bits_size,
	auto_buffer_in_a_bits_source,
	auto_buffer_in_a_bits_address,
	auto_buffer_in_a_bits_mask,
	auto_buffer_in_a_bits_corrupt,
	auto_buffer_in_d_ready,
	auto_buffer_in_d_valid,
	auto_buffer_in_d_bits_opcode,
	auto_buffer_in_d_bits_param,
	auto_buffer_in_d_bits_size,
	auto_buffer_in_d_bits_source,
	auto_buffer_in_d_bits_sink,
	auto_buffer_in_d_bits_denied,
	auto_buffer_in_d_bits_data,
	auto_buffer_in_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_buffer_in_a_ready;
	input auto_buffer_in_a_valid;
	input [2:0] auto_buffer_in_a_bits_opcode;
	input [2:0] auto_buffer_in_a_bits_param;
	input [3:0] auto_buffer_in_a_bits_size;
	input [2:0] auto_buffer_in_a_bits_source;
	input [13:0] auto_buffer_in_a_bits_address;
	input [3:0] auto_buffer_in_a_bits_mask;
	input auto_buffer_in_a_bits_corrupt;
	input auto_buffer_in_d_ready;
	output wire auto_buffer_in_d_valid;
	output wire [2:0] auto_buffer_in_d_bits_opcode;
	output wire [1:0] auto_buffer_in_d_bits_param;
	output wire [3:0] auto_buffer_in_d_bits_size;
	output wire [2:0] auto_buffer_in_d_bits_source;
	output wire auto_buffer_in_d_bits_sink;
	output wire auto_buffer_in_d_bits_denied;
	output wire [31:0] auto_buffer_in_d_bits_data;
	output wire auto_buffer_in_d_bits_corrupt;
	wire error_clock;
	wire error_reset;
	wire error_auto_in_a_ready;
	wire error_auto_in_a_valid;
	wire [2:0] error_auto_in_a_bits_opcode;
	wire [2:0] error_auto_in_a_bits_param;
	wire [3:0] error_auto_in_a_bits_size;
	wire [2:0] error_auto_in_a_bits_source;
	wire [13:0] error_auto_in_a_bits_address;
	wire [3:0] error_auto_in_a_bits_mask;
	wire error_auto_in_a_bits_corrupt;
	wire error_auto_in_d_ready;
	wire error_auto_in_d_valid;
	wire [2:0] error_auto_in_d_bits_opcode;
	wire [3:0] error_auto_in_d_bits_size;
	wire [2:0] error_auto_in_d_bits_source;
	wire error_auto_in_d_bits_corrupt;
	wire buffer_clock;
	wire buffer_reset;
	wire buffer_auto_in_a_ready;
	wire buffer_auto_in_a_valid;
	wire [2:0] buffer_auto_in_a_bits_opcode;
	wire [2:0] buffer_auto_in_a_bits_param;
	wire [3:0] buffer_auto_in_a_bits_size;
	wire [2:0] buffer_auto_in_a_bits_source;
	wire [13:0] buffer_auto_in_a_bits_address;
	wire [3:0] buffer_auto_in_a_bits_mask;
	wire buffer_auto_in_a_bits_corrupt;
	wire buffer_auto_in_d_ready;
	wire buffer_auto_in_d_valid;
	wire [2:0] buffer_auto_in_d_bits_opcode;
	wire [1:0] buffer_auto_in_d_bits_param;
	wire [3:0] buffer_auto_in_d_bits_size;
	wire [2:0] buffer_auto_in_d_bits_source;
	wire buffer_auto_in_d_bits_sink;
	wire buffer_auto_in_d_bits_denied;
	wire [31:0] buffer_auto_in_d_bits_data;
	wire buffer_auto_in_d_bits_corrupt;
	wire buffer_auto_out_a_ready;
	wire buffer_auto_out_a_valid;
	wire [2:0] buffer_auto_out_a_bits_opcode;
	wire [2:0] buffer_auto_out_a_bits_param;
	wire [3:0] buffer_auto_out_a_bits_size;
	wire [2:0] buffer_auto_out_a_bits_source;
	wire [13:0] buffer_auto_out_a_bits_address;
	wire [3:0] buffer_auto_out_a_bits_mask;
	wire buffer_auto_out_a_bits_corrupt;
	wire buffer_auto_out_d_ready;
	wire buffer_auto_out_d_valid;
	wire [2:0] buffer_auto_out_d_bits_opcode;
	wire [3:0] buffer_auto_out_d_bits_size;
	wire [2:0] buffer_auto_out_d_bits_source;
	wire buffer_auto_out_d_bits_corrupt;
	TLError error(
		.clock(error_clock),
		.reset(error_reset),
		.auto_in_a_ready(error_auto_in_a_ready),
		.auto_in_a_valid(error_auto_in_a_valid),
		.auto_in_a_bits_opcode(error_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(error_auto_in_a_bits_param),
		.auto_in_a_bits_size(error_auto_in_a_bits_size),
		.auto_in_a_bits_source(error_auto_in_a_bits_source),
		.auto_in_a_bits_address(error_auto_in_a_bits_address),
		.auto_in_a_bits_mask(error_auto_in_a_bits_mask),
		.auto_in_a_bits_corrupt(error_auto_in_a_bits_corrupt),
		.auto_in_d_ready(error_auto_in_d_ready),
		.auto_in_d_valid(error_auto_in_d_valid),
		.auto_in_d_bits_opcode(error_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(error_auto_in_d_bits_size),
		.auto_in_d_bits_source(error_auto_in_d_bits_source),
		.auto_in_d_bits_corrupt(error_auto_in_d_bits_corrupt)
	);
	TLBuffer_7 buffer(
		.clock(buffer_clock),
		.reset(buffer_reset),
		.auto_in_a_ready(buffer_auto_in_a_ready),
		.auto_in_a_valid(buffer_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
		.auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_auto_in_d_ready),
		.auto_in_d_valid(buffer_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_auto_out_a_ready),
		.auto_out_a_valid(buffer_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
		.auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_auto_out_d_ready),
		.auto_out_d_valid(buffer_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(buffer_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_auto_out_d_bits_source),
		.auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt)
	);
	assign auto_buffer_in_a_ready = buffer_auto_in_a_ready;
	assign auto_buffer_in_d_valid = buffer_auto_in_d_valid;
	assign auto_buffer_in_d_bits_opcode = buffer_auto_in_d_bits_opcode;
	assign auto_buffer_in_d_bits_param = buffer_auto_in_d_bits_param;
	assign auto_buffer_in_d_bits_size = buffer_auto_in_d_bits_size;
	assign auto_buffer_in_d_bits_source = buffer_auto_in_d_bits_source;
	assign auto_buffer_in_d_bits_sink = buffer_auto_in_d_bits_sink;
	assign auto_buffer_in_d_bits_denied = buffer_auto_in_d_bits_denied;
	assign auto_buffer_in_d_bits_data = buffer_auto_in_d_bits_data;
	assign auto_buffer_in_d_bits_corrupt = buffer_auto_in_d_bits_corrupt;
	assign error_clock = clock;
	assign error_reset = reset;
	assign error_auto_in_a_valid = buffer_auto_out_a_valid;
	assign error_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode;
	assign error_auto_in_a_bits_param = buffer_auto_out_a_bits_param;
	assign error_auto_in_a_bits_size = buffer_auto_out_a_bits_size;
	assign error_auto_in_a_bits_source = buffer_auto_out_a_bits_source;
	assign error_auto_in_a_bits_address = buffer_auto_out_a_bits_address;
	assign error_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask;
	assign error_auto_in_a_bits_corrupt = buffer_auto_out_a_bits_corrupt;
	assign error_auto_in_d_ready = buffer_auto_out_d_ready;
	assign buffer_clock = clock;
	assign buffer_reset = reset;
	assign buffer_auto_in_a_valid = auto_buffer_in_a_valid;
	assign buffer_auto_in_a_bits_opcode = auto_buffer_in_a_bits_opcode;
	assign buffer_auto_in_a_bits_param = auto_buffer_in_a_bits_param;
	assign buffer_auto_in_a_bits_size = auto_buffer_in_a_bits_size;
	assign buffer_auto_in_a_bits_source = auto_buffer_in_a_bits_source;
	assign buffer_auto_in_a_bits_address = auto_buffer_in_a_bits_address;
	assign buffer_auto_in_a_bits_mask = auto_buffer_in_a_bits_mask;
	assign buffer_auto_in_a_bits_corrupt = auto_buffer_in_a_bits_corrupt;
	assign buffer_auto_in_d_ready = auto_buffer_in_d_ready;
	assign buffer_auto_out_a_ready = error_auto_in_a_ready;
	assign buffer_auto_out_d_valid = error_auto_in_d_valid;
	assign buffer_auto_out_d_bits_opcode = error_auto_in_d_bits_opcode;
	assign buffer_auto_out_d_bits_size = error_auto_in_d_bits_size;
	assign buffer_auto_out_d_bits_source = error_auto_in_d_bits_source;
	assign buffer_auto_out_d_bits_corrupt = error_auto_in_d_bits_corrupt;
endmodule
module TLBuffer_8 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input [1:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire [1:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire [1:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input [1:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module TLWidthWidget_5 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [30:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [30:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module TLInterconnectCoupler_9 (
	auto_widget_in_a_ready,
	auto_widget_in_a_valid,
	auto_widget_in_a_bits_opcode,
	auto_widget_in_a_bits_param,
	auto_widget_in_a_bits_size,
	auto_widget_in_a_bits_source,
	auto_widget_in_a_bits_address,
	auto_widget_in_a_bits_mask,
	auto_widget_in_a_bits_data,
	auto_widget_in_a_bits_corrupt,
	auto_widget_in_d_ready,
	auto_widget_in_d_valid,
	auto_widget_in_d_bits_opcode,
	auto_widget_in_d_bits_param,
	auto_widget_in_d_bits_size,
	auto_widget_in_d_bits_source,
	auto_widget_in_d_bits_sink,
	auto_widget_in_d_bits_denied,
	auto_widget_in_d_bits_data,
	auto_widget_in_d_bits_corrupt,
	auto_bus_xing_out_a_ready,
	auto_bus_xing_out_a_valid,
	auto_bus_xing_out_a_bits_opcode,
	auto_bus_xing_out_a_bits_param,
	auto_bus_xing_out_a_bits_size,
	auto_bus_xing_out_a_bits_source,
	auto_bus_xing_out_a_bits_address,
	auto_bus_xing_out_a_bits_mask,
	auto_bus_xing_out_a_bits_data,
	auto_bus_xing_out_a_bits_corrupt,
	auto_bus_xing_out_d_ready,
	auto_bus_xing_out_d_valid,
	auto_bus_xing_out_d_bits_opcode,
	auto_bus_xing_out_d_bits_param,
	auto_bus_xing_out_d_bits_size,
	auto_bus_xing_out_d_bits_source,
	auto_bus_xing_out_d_bits_sink,
	auto_bus_xing_out_d_bits_denied,
	auto_bus_xing_out_d_bits_data,
	auto_bus_xing_out_d_bits_corrupt
);
	output wire auto_widget_in_a_ready;
	input auto_widget_in_a_valid;
	input [2:0] auto_widget_in_a_bits_opcode;
	input [2:0] auto_widget_in_a_bits_param;
	input [2:0] auto_widget_in_a_bits_size;
	input [2:0] auto_widget_in_a_bits_source;
	input [30:0] auto_widget_in_a_bits_address;
	input [3:0] auto_widget_in_a_bits_mask;
	input [31:0] auto_widget_in_a_bits_data;
	input auto_widget_in_a_bits_corrupt;
	input auto_widget_in_d_ready;
	output wire auto_widget_in_d_valid;
	output wire [2:0] auto_widget_in_d_bits_opcode;
	output wire [1:0] auto_widget_in_d_bits_param;
	output wire [2:0] auto_widget_in_d_bits_size;
	output wire [2:0] auto_widget_in_d_bits_source;
	output wire auto_widget_in_d_bits_sink;
	output wire auto_widget_in_d_bits_denied;
	output wire [31:0] auto_widget_in_d_bits_data;
	output wire auto_widget_in_d_bits_corrupt;
	input auto_bus_xing_out_a_ready;
	output wire auto_bus_xing_out_a_valid;
	output wire [2:0] auto_bus_xing_out_a_bits_opcode;
	output wire [2:0] auto_bus_xing_out_a_bits_param;
	output wire [2:0] auto_bus_xing_out_a_bits_size;
	output wire [2:0] auto_bus_xing_out_a_bits_source;
	output wire [30:0] auto_bus_xing_out_a_bits_address;
	output wire [3:0] auto_bus_xing_out_a_bits_mask;
	output wire [31:0] auto_bus_xing_out_a_bits_data;
	output wire auto_bus_xing_out_a_bits_corrupt;
	output wire auto_bus_xing_out_d_ready;
	input auto_bus_xing_out_d_valid;
	input [2:0] auto_bus_xing_out_d_bits_opcode;
	input [1:0] auto_bus_xing_out_d_bits_param;
	input [2:0] auto_bus_xing_out_d_bits_size;
	input [2:0] auto_bus_xing_out_d_bits_source;
	input auto_bus_xing_out_d_bits_sink;
	input auto_bus_xing_out_d_bits_denied;
	input [31:0] auto_bus_xing_out_d_bits_data;
	input auto_bus_xing_out_d_bits_corrupt;
	wire widget_auto_in_a_ready;
	wire widget_auto_in_a_valid;
	wire [2:0] widget_auto_in_a_bits_opcode;
	wire [2:0] widget_auto_in_a_bits_param;
	wire [2:0] widget_auto_in_a_bits_size;
	wire [2:0] widget_auto_in_a_bits_source;
	wire [30:0] widget_auto_in_a_bits_address;
	wire [3:0] widget_auto_in_a_bits_mask;
	wire [31:0] widget_auto_in_a_bits_data;
	wire widget_auto_in_a_bits_corrupt;
	wire widget_auto_in_d_ready;
	wire widget_auto_in_d_valid;
	wire [2:0] widget_auto_in_d_bits_opcode;
	wire [1:0] widget_auto_in_d_bits_param;
	wire [2:0] widget_auto_in_d_bits_size;
	wire [2:0] widget_auto_in_d_bits_source;
	wire widget_auto_in_d_bits_sink;
	wire widget_auto_in_d_bits_denied;
	wire [31:0] widget_auto_in_d_bits_data;
	wire widget_auto_in_d_bits_corrupt;
	wire widget_auto_out_a_ready;
	wire widget_auto_out_a_valid;
	wire [2:0] widget_auto_out_a_bits_opcode;
	wire [2:0] widget_auto_out_a_bits_param;
	wire [2:0] widget_auto_out_a_bits_size;
	wire [2:0] widget_auto_out_a_bits_source;
	wire [30:0] widget_auto_out_a_bits_address;
	wire [3:0] widget_auto_out_a_bits_mask;
	wire [31:0] widget_auto_out_a_bits_data;
	wire widget_auto_out_a_bits_corrupt;
	wire widget_auto_out_d_ready;
	wire widget_auto_out_d_valid;
	wire [2:0] widget_auto_out_d_bits_opcode;
	wire [1:0] widget_auto_out_d_bits_param;
	wire [2:0] widget_auto_out_d_bits_size;
	wire [2:0] widget_auto_out_d_bits_source;
	wire widget_auto_out_d_bits_sink;
	wire widget_auto_out_d_bits_denied;
	wire [31:0] widget_auto_out_d_bits_data;
	wire widget_auto_out_d_bits_corrupt;
	TLWidthWidget_5 widget(
		.auto_in_a_ready(widget_auto_in_a_ready),
		.auto_in_a_valid(widget_auto_in_a_valid),
		.auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(widget_auto_in_a_bits_param),
		.auto_in_a_bits_size(widget_auto_in_a_bits_size),
		.auto_in_a_bits_source(widget_auto_in_a_bits_source),
		.auto_in_a_bits_address(widget_auto_in_a_bits_address),
		.auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
		.auto_in_a_bits_data(widget_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(widget_auto_in_a_bits_corrupt),
		.auto_in_d_ready(widget_auto_in_d_ready),
		.auto_in_d_valid(widget_auto_in_d_valid),
		.auto_in_d_bits_opcode(widget_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(widget_auto_in_d_bits_param),
		.auto_in_d_bits_size(widget_auto_in_d_bits_size),
		.auto_in_d_bits_source(widget_auto_in_d_bits_source),
		.auto_in_d_bits_sink(widget_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(widget_auto_in_d_bits_denied),
		.auto_in_d_bits_data(widget_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(widget_auto_in_d_bits_corrupt),
		.auto_out_a_ready(widget_auto_out_a_ready),
		.auto_out_a_valid(widget_auto_out_a_valid),
		.auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(widget_auto_out_a_bits_param),
		.auto_out_a_bits_size(widget_auto_out_a_bits_size),
		.auto_out_a_bits_source(widget_auto_out_a_bits_source),
		.auto_out_a_bits_address(widget_auto_out_a_bits_address),
		.auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
		.auto_out_a_bits_data(widget_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(widget_auto_out_a_bits_corrupt),
		.auto_out_d_ready(widget_auto_out_d_ready),
		.auto_out_d_valid(widget_auto_out_d_valid),
		.auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(widget_auto_out_d_bits_param),
		.auto_out_d_bits_size(widget_auto_out_d_bits_size),
		.auto_out_d_bits_source(widget_auto_out_d_bits_source),
		.auto_out_d_bits_sink(widget_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(widget_auto_out_d_bits_denied),
		.auto_out_d_bits_data(widget_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(widget_auto_out_d_bits_corrupt)
	);
	assign auto_widget_in_a_ready = widget_auto_in_a_ready;
	assign auto_widget_in_d_valid = widget_auto_in_d_valid;
	assign auto_widget_in_d_bits_opcode = widget_auto_in_d_bits_opcode;
	assign auto_widget_in_d_bits_param = widget_auto_in_d_bits_param;
	assign auto_widget_in_d_bits_size = widget_auto_in_d_bits_size;
	assign auto_widget_in_d_bits_source = widget_auto_in_d_bits_source;
	assign auto_widget_in_d_bits_sink = widget_auto_in_d_bits_sink;
	assign auto_widget_in_d_bits_denied = widget_auto_in_d_bits_denied;
	assign auto_widget_in_d_bits_data = widget_auto_in_d_bits_data;
	assign auto_widget_in_d_bits_corrupt = widget_auto_in_d_bits_corrupt;
	assign auto_bus_xing_out_a_valid = widget_auto_out_a_valid;
	assign auto_bus_xing_out_a_bits_opcode = widget_auto_out_a_bits_opcode;
	assign auto_bus_xing_out_a_bits_param = widget_auto_out_a_bits_param;
	assign auto_bus_xing_out_a_bits_size = widget_auto_out_a_bits_size;
	assign auto_bus_xing_out_a_bits_source = widget_auto_out_a_bits_source;
	assign auto_bus_xing_out_a_bits_address = widget_auto_out_a_bits_address;
	assign auto_bus_xing_out_a_bits_mask = widget_auto_out_a_bits_mask;
	assign auto_bus_xing_out_a_bits_data = widget_auto_out_a_bits_data;
	assign auto_bus_xing_out_a_bits_corrupt = widget_auto_out_a_bits_corrupt;
	assign auto_bus_xing_out_d_ready = widget_auto_out_d_ready;
	assign widget_auto_in_a_valid = auto_widget_in_a_valid;
	assign widget_auto_in_a_bits_opcode = auto_widget_in_a_bits_opcode;
	assign widget_auto_in_a_bits_param = auto_widget_in_a_bits_param;
	assign widget_auto_in_a_bits_size = auto_widget_in_a_bits_size;
	assign widget_auto_in_a_bits_source = auto_widget_in_a_bits_source;
	assign widget_auto_in_a_bits_address = auto_widget_in_a_bits_address;
	assign widget_auto_in_a_bits_mask = auto_widget_in_a_bits_mask;
	assign widget_auto_in_a_bits_data = auto_widget_in_a_bits_data;
	assign widget_auto_in_a_bits_corrupt = auto_widget_in_a_bits_corrupt;
	assign widget_auto_in_d_ready = auto_widget_in_d_ready;
	assign widget_auto_out_a_ready = auto_bus_xing_out_a_ready;
	assign widget_auto_out_d_valid = auto_bus_xing_out_d_valid;
	assign widget_auto_out_d_bits_opcode = auto_bus_xing_out_d_bits_opcode;
	assign widget_auto_out_d_bits_param = auto_bus_xing_out_d_bits_param;
	assign widget_auto_out_d_bits_size = auto_bus_xing_out_d_bits_size;
	assign widget_auto_out_d_bits_source = auto_bus_xing_out_d_bits_source;
	assign widget_auto_out_d_bits_sink = auto_bus_xing_out_d_bits_sink;
	assign widget_auto_out_d_bits_denied = auto_bus_xing_out_d_bits_denied;
	assign widget_auto_out_d_bits_data = auto_bus_xing_out_d_bits_data;
	assign widget_auto_out_d_bits_corrupt = auto_bus_xing_out_d_bits_corrupt;
endmodule
module TLMonitor_23 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [27:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [27:0] _GEN_71 = {22'd0, is_aligned_mask};
	wire [27:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 28'h0000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [27:0] _T_56 = io_in_a_bits_address ^ 28'hc000000;
	wire [28:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [28:0] _T_59 = $signed(_T_57) & -29'sh04000000;
	wire _T_60 = $signed(_T_59) == 29'sh00000000;
	wire _T_92 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_96 = ~io_in_a_bits_mask;
	wire _T_97 = _T_96 == 4'h0;
	wire _T_101 = ~io_in_a_bits_corrupt;
	wire _T_105 = io_in_a_bits_opcode == 3'h7;
	wire _T_159 = io_in_a_bits_param != 3'h0;
	wire _T_172 = io_in_a_bits_opcode == 3'h4;
	wire _T_189 = io_in_a_bits_size <= 3'h6;
	wire _T_197 = _T_189 & _T_60;
	wire _T_208 = io_in_a_bits_param == 3'h0;
	wire _T_212 = io_in_a_bits_mask == mask;
	wire _T_220 = io_in_a_bits_opcode == 3'h0;
	wire _T_244 = source_ok & _T_197;
	wire _T_262 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_300 = ~mask;
	wire [3:0] _T_301 = io_in_a_bits_mask & _T_300;
	wire _T_302 = _T_301 == 4'h0;
	wire _T_306 = io_in_a_bits_opcode == 3'h2;
	wire _T_337 = io_in_a_bits_param <= 3'h4;
	wire _T_345 = io_in_a_bits_opcode == 3'h3;
	wire _T_376 = io_in_a_bits_param <= 3'h3;
	wire _T_384 = io_in_a_bits_opcode == 3'h5;
	wire _T_415 = io_in_a_bits_param <= 3'h1;
	wire _T_427 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_431 = io_in_d_bits_opcode == 3'h6;
	wire _T_435 = io_in_d_bits_size >= 3'h2;
	wire _T_451 = io_in_d_bits_opcode == 3'h4;
	wire _T_479 = io_in_d_bits_opcode == 3'h5;
	wire _T_508 = io_in_d_bits_opcode == 3'h0;
	wire _T_525 = io_in_d_bits_opcode == 3'h1;
	wire _T_543 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [27:0] address;
	wire _T_573 = io_in_a_valid & ~a_first;
	wire _T_574 = io_in_a_bits_opcode == opcode;
	wire _T_578 = io_in_a_bits_param == param;
	wire _T_582 = io_in_a_bits_size == size;
	wire _T_586 = io_in_a_bits_source == source;
	wire _T_590 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	wire _T_597 = io_in_d_valid & ~d_first;
	wire _T_598 = io_in_d_bits_opcode == opcode_1;
	wire _T_606 = io_in_d_bits_size == size_1;
	wire _T_610 = io_in_d_bits_source == source_1;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_624 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire [7:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire _T_627 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_629 = inflight >> io_in_a_bits_source;
	wire _T_631 = ~_T_629[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_635 = io_in_d_valid & d_first_1;
	wire _T_637 = ~_T_431;
	wire _T_638 = (io_in_d_valid & d_first_1) & ~_T_431;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [7:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_431 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_637 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_637 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_624 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_648 = inflight >> io_in_d_bits_source;
	wire _T_650 = _T_648[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_655 = io_in_d_bits_opcode == _GEN_40;
	wire _T_656 = (io_in_d_bits_opcode == _GEN_32) | _T_655;
	wire _T_660 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_667 = io_in_d_bits_opcode == _GEN_56;
	wire _T_668 = (io_in_d_bits_opcode == _GEN_48) | _T_667;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_672 = _GEN_82 == a_size_lookup;
	wire _T_682 = (((_T_635 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_637;
	wire _T_684 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set_wo_ready = _GEN_15[4:0];
	wire [4:0] d_clr_wo_ready = _GEN_21[4:0];
	wire _T_691 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_700 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_726 = (io_in_d_valid & d_first_2) & _T_431;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_431 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_431 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_734 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_744 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_769 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Repeater_3 (
	clock,
	reset,
	io_repeat,
	io_full,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	input io_repeat;
	output wire io_full;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [27:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [27:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire io_deq_bits_corrupt;
	reg full;
	reg [2:0] saved_opcode;
	reg [2:0] saved_param;
	reg [2:0] saved_size;
	reg [2:0] saved_source;
	reg [27:0] saved_address;
	reg [3:0] saved_mask;
	reg saved_corrupt;
	wire _T = io_enq_ready & io_enq_valid;
	wire _GEN_0 = (_T & io_repeat) | full;
	wire _T_2 = io_deq_ready & io_deq_valid;
	assign io_full = full;
	assign io_enq_ready = io_deq_ready & ~full;
	assign io_deq_valid = io_enq_valid | full;
	assign io_deq_bits_opcode = (full ? saved_opcode : io_enq_bits_opcode);
	assign io_deq_bits_param = (full ? saved_param : io_enq_bits_param);
	assign io_deq_bits_size = (full ? saved_size : io_enq_bits_size);
	assign io_deq_bits_source = (full ? saved_source : io_enq_bits_source);
	assign io_deq_bits_address = (full ? saved_address : io_enq_bits_address);
	assign io_deq_bits_mask = (full ? saved_mask : io_enq_bits_mask);
	assign io_deq_bits_corrupt = (full ? saved_corrupt : io_enq_bits_corrupt);
	always @(posedge clock) begin
		if (reset)
			full <= 1'h0;
		else if (_T_2 & ~io_repeat)
			full <= 1'h0;
		else
			full <= _GEN_0;
		if (_T & io_repeat)
			saved_opcode <= io_enq_bits_opcode;
		if (_T & io_repeat)
			saved_param <= io_enq_bits_param;
		if (_T & io_repeat)
			saved_size <= io_enq_bits_size;
		if (_T & io_repeat)
			saved_source <= io_enq_bits_source;
		if (_T & io_repeat)
			saved_address <= io_enq_bits_address;
		if (_T & io_repeat)
			saved_mask <= io_enq_bits_mask;
		if (_T & io_repeat)
			saved_corrupt <= io_enq_bits_corrupt;
	end
endmodule
module TLFragmenter_2 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [27:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire [7:0] auto_out_a_bits_source;
	output wire [27:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_size;
	input [7:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [27:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire repeater_clock;
	wire repeater_reset;
	wire repeater_io_repeat;
	wire repeater_io_full;
	wire repeater_io_enq_ready;
	wire repeater_io_enq_valid;
	wire [2:0] repeater_io_enq_bits_opcode;
	wire [2:0] repeater_io_enq_bits_param;
	wire [2:0] repeater_io_enq_bits_size;
	wire [2:0] repeater_io_enq_bits_source;
	wire [27:0] repeater_io_enq_bits_address;
	wire [3:0] repeater_io_enq_bits_mask;
	wire repeater_io_enq_bits_corrupt;
	wire repeater_io_deq_ready;
	wire repeater_io_deq_valid;
	wire [2:0] repeater_io_deq_bits_opcode;
	wire [2:0] repeater_io_deq_bits_param;
	wire [2:0] repeater_io_deq_bits_size;
	wire [2:0] repeater_io_deq_bits_source;
	wire [27:0] repeater_io_deq_bits_address;
	wire [3:0] repeater_io_deq_bits_mask;
	wire repeater_io_deq_bits_corrupt;
	reg [3:0] acknum;
	reg [2:0] dOrig;
	reg dToggle;
	wire [3:0] dFragnum = auto_out_d_bits_source[3:0];
	wire dFirst = acknum == 4'h0;
	wire dLast = dFragnum == 4'h0;
	wire [3:0] _dsizeOH_T = 4'h1 << auto_out_d_bits_size;
	wire [2:0] dsizeOH = _dsizeOH_T[2:0];
	wire [4:0] _dsizeOH1_T_1 = 5'h03 << auto_out_d_bits_size;
	wire [1:0] dsizeOH1 = ~_dsizeOH1_T_1[1:0];
	wire dHasData = auto_out_d_bits_opcode[0];
	wire _T_5 = ~reset;
	wire ack_decrement = dHasData | dsizeOH[2];
	wire [5:0] _dFirst_size_T = {dFragnum, 2'h0};
	wire [5:0] _GEN_7 = {4'd0, dsizeOH1};
	wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7;
	wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0};
	wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h01;
	wire [6:0] _dFirst_size_T_4 = {1'h0, _dFirst_size_T_1};
	wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4;
	wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5;
	wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4];
	wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0];
	wire _dFirst_size_T_7 = |dFirst_size_hi;
	wire [3:0] _GEN_8 = {1'd0, dFirst_size_hi};
	wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo;
	wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2];
	wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0];
	wire _dFirst_size_T_9 = |dFirst_size_hi_1;
	wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1;
	wire [2:0] dFirst_size = {_dFirst_size_T_7, _dFirst_size_T_9, _dFirst_size_T_10[1]};
	wire drop = ~dHasData & ~dLast;
	wire bundleOut_0_d_ready = auto_in_d_ready | drop;
	wire _T_7 = bundleOut_0_d_ready & auto_out_d_valid;
	wire [3:0] _GEN_9 = {3'd0, ack_decrement};
	wire [3:0] _acknum_T_1 = acknum - _GEN_9;
	wire [2:0] aFrag = (repeater_io_deq_bits_size > 3'h2 ? 3'h2 : repeater_io_deq_bits_size);
	wire [12:0] _aOrigOH1_T_1 = 13'h003f << repeater_io_deq_bits_size;
	wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0];
	wire [8:0] _aFragOH1_T_1 = 9'h003 << aFrag;
	wire [1:0] aFragOH1 = ~_aFragOH1_T_1[1:0];
	wire aHasData = ~repeater_io_deq_bits_opcode[2];
	reg [3:0] gennum;
	wire aFirst = gennum == 4'h0;
	wire [3:0] _old_gennum1_T_2 = gennum - 4'h1;
	wire [3:0] old_gennum1 = (aFirst ? aOrigOH1[5:2] : _old_gennum1_T_2);
	wire [3:0] _new_gennum_T = ~old_gennum1;
	wire [3:0] new_gennum = ~_new_gennum_T;
	reg aToggle_r;
	wire _GEN_5 = (aFirst ? dToggle : aToggle_r);
	wire aToggle = ~_GEN_5;
	wire bundleOut_0_a_valid = repeater_io_deq_valid;
	wire _T_8 = auto_out_a_ready & bundleOut_0_a_valid;
	wire _repeater_io_repeat_T = ~aHasData;
	wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 2'h0};
	wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1;
	wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1;
	wire [5:0] _GEN_10 = {4'd0, aFragOH1};
	wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10;
	wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h03;
	wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4;
	wire [27:0] _GEN_11 = {22'd0, _bundleOut_0_a_bits_address_T_5};
	wire [3:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source, aToggle};
	wire _T_9 = ~repeater_io_full;
	TLMonitor_23 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	Repeater_3 repeater(
		.clock(repeater_clock),
		.reset(repeater_reset),
		.io_repeat(repeater_io_repeat),
		.io_full(repeater_io_full),
		.io_enq_ready(repeater_io_enq_ready),
		.io_enq_valid(repeater_io_enq_valid),
		.io_enq_bits_opcode(repeater_io_enq_bits_opcode),
		.io_enq_bits_param(repeater_io_enq_bits_param),
		.io_enq_bits_size(repeater_io_enq_bits_size),
		.io_enq_bits_source(repeater_io_enq_bits_source),
		.io_enq_bits_address(repeater_io_enq_bits_address),
		.io_enq_bits_mask(repeater_io_enq_bits_mask),
		.io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
		.io_deq_ready(repeater_io_deq_ready),
		.io_deq_valid(repeater_io_deq_valid),
		.io_deq_bits_opcode(repeater_io_deq_bits_opcode),
		.io_deq_bits_param(repeater_io_deq_bits_param),
		.io_deq_bits_size(repeater_io_deq_bits_size),
		.io_deq_bits_source(repeater_io_deq_bits_source),
		.io_deq_bits_address(repeater_io_deq_bits_address),
		.io_deq_bits_mask(repeater_io_deq_bits_mask),
		.io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = repeater_io_enq_ready;
	assign auto_in_d_valid = auto_out_d_valid & ~drop;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign auto_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_out_a_valid = repeater_io_deq_valid;
	assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode;
	assign auto_out_a_bits_param = repeater_io_deq_bits_param;
	assign auto_out_a_bits_size = aFrag[1:0];
	assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi, new_gennum};
	assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11;
	assign auto_out_a_bits_mask = (repeater_io_full ? 4'hf : auto_in_a_bits_mask);
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready | drop;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = repeater_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid & ~drop;
	assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_io_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign repeater_clock = clock;
	assign repeater_reset = reset;
	assign repeater_io_repeat = ~aHasData & (new_gennum != 4'h0);
	assign repeater_io_enq_valid = auto_in_a_valid;
	assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign repeater_io_enq_bits_param = auto_in_a_bits_param;
	assign repeater_io_enq_bits_size = auto_in_a_bits_size;
	assign repeater_io_enq_bits_source = auto_in_a_bits_source;
	assign repeater_io_enq_bits_address = auto_in_a_bits_address;
	assign repeater_io_enq_bits_mask = auto_in_a_bits_mask;
	assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign repeater_io_deq_ready = auto_out_a_ready;
	always @(posedge clock) begin
		if (reset)
			acknum <= 4'h0;
		else if (_T_7)
			if (dFirst)
				acknum <= dFragnum;
			else
				acknum <= _acknum_T_1;
		if (_T_7)
			if (dFirst)
				dOrig <= dFirst_size;
		if (reset)
			dToggle <= 1'h0;
		else if (_T_7)
			if (dFirst)
				dToggle <= auto_out_d_bits_source[4];
		if (reset)
			gennum <= 4'h0;
		else if (_T_8)
			gennum <= new_gennum;
		if (aFirst)
			aToggle_r <= dToggle;
	end
endmodule
module TLInterconnectCoupler_10 (
	clock,
	reset,
	auto_fragmenter_out_a_ready,
	auto_fragmenter_out_a_valid,
	auto_fragmenter_out_a_bits_opcode,
	auto_fragmenter_out_a_bits_param,
	auto_fragmenter_out_a_bits_size,
	auto_fragmenter_out_a_bits_source,
	auto_fragmenter_out_a_bits_address,
	auto_fragmenter_out_a_bits_mask,
	auto_fragmenter_out_a_bits_data,
	auto_fragmenter_out_a_bits_corrupt,
	auto_fragmenter_out_d_ready,
	auto_fragmenter_out_d_valid,
	auto_fragmenter_out_d_bits_opcode,
	auto_fragmenter_out_d_bits_size,
	auto_fragmenter_out_d_bits_source,
	auto_fragmenter_out_d_bits_data,
	auto_tl_in_a_ready,
	auto_tl_in_a_valid,
	auto_tl_in_a_bits_opcode,
	auto_tl_in_a_bits_param,
	auto_tl_in_a_bits_size,
	auto_tl_in_a_bits_source,
	auto_tl_in_a_bits_address,
	auto_tl_in_a_bits_mask,
	auto_tl_in_a_bits_data,
	auto_tl_in_a_bits_corrupt,
	auto_tl_in_d_ready,
	auto_tl_in_d_valid,
	auto_tl_in_d_bits_opcode,
	auto_tl_in_d_bits_size,
	auto_tl_in_d_bits_source,
	auto_tl_in_d_bits_data
);
	input clock;
	input reset;
	input auto_fragmenter_out_a_ready;
	output wire auto_fragmenter_out_a_valid;
	output wire [2:0] auto_fragmenter_out_a_bits_opcode;
	output wire [2:0] auto_fragmenter_out_a_bits_param;
	output wire [1:0] auto_fragmenter_out_a_bits_size;
	output wire [7:0] auto_fragmenter_out_a_bits_source;
	output wire [27:0] auto_fragmenter_out_a_bits_address;
	output wire [3:0] auto_fragmenter_out_a_bits_mask;
	output wire [31:0] auto_fragmenter_out_a_bits_data;
	output wire auto_fragmenter_out_a_bits_corrupt;
	output wire auto_fragmenter_out_d_ready;
	input auto_fragmenter_out_d_valid;
	input [2:0] auto_fragmenter_out_d_bits_opcode;
	input [1:0] auto_fragmenter_out_d_bits_size;
	input [7:0] auto_fragmenter_out_d_bits_source;
	input [31:0] auto_fragmenter_out_d_bits_data;
	output wire auto_tl_in_a_ready;
	input auto_tl_in_a_valid;
	input [2:0] auto_tl_in_a_bits_opcode;
	input [2:0] auto_tl_in_a_bits_param;
	input [2:0] auto_tl_in_a_bits_size;
	input [2:0] auto_tl_in_a_bits_source;
	input [27:0] auto_tl_in_a_bits_address;
	input [3:0] auto_tl_in_a_bits_mask;
	input [31:0] auto_tl_in_a_bits_data;
	input auto_tl_in_a_bits_corrupt;
	input auto_tl_in_d_ready;
	output wire auto_tl_in_d_valid;
	output wire [2:0] auto_tl_in_d_bits_opcode;
	output wire [2:0] auto_tl_in_d_bits_size;
	output wire [2:0] auto_tl_in_d_bits_source;
	output wire [31:0] auto_tl_in_d_bits_data;
	wire fragmenter_clock;
	wire fragmenter_reset;
	wire fragmenter_auto_in_a_ready;
	wire fragmenter_auto_in_a_valid;
	wire [2:0] fragmenter_auto_in_a_bits_opcode;
	wire [2:0] fragmenter_auto_in_a_bits_param;
	wire [2:0] fragmenter_auto_in_a_bits_size;
	wire [2:0] fragmenter_auto_in_a_bits_source;
	wire [27:0] fragmenter_auto_in_a_bits_address;
	wire [3:0] fragmenter_auto_in_a_bits_mask;
	wire [31:0] fragmenter_auto_in_a_bits_data;
	wire fragmenter_auto_in_a_bits_corrupt;
	wire fragmenter_auto_in_d_ready;
	wire fragmenter_auto_in_d_valid;
	wire [2:0] fragmenter_auto_in_d_bits_opcode;
	wire [2:0] fragmenter_auto_in_d_bits_size;
	wire [2:0] fragmenter_auto_in_d_bits_source;
	wire [31:0] fragmenter_auto_in_d_bits_data;
	wire fragmenter_auto_out_a_ready;
	wire fragmenter_auto_out_a_valid;
	wire [2:0] fragmenter_auto_out_a_bits_opcode;
	wire [2:0] fragmenter_auto_out_a_bits_param;
	wire [1:0] fragmenter_auto_out_a_bits_size;
	wire [7:0] fragmenter_auto_out_a_bits_source;
	wire [27:0] fragmenter_auto_out_a_bits_address;
	wire [3:0] fragmenter_auto_out_a_bits_mask;
	wire [31:0] fragmenter_auto_out_a_bits_data;
	wire fragmenter_auto_out_a_bits_corrupt;
	wire fragmenter_auto_out_d_ready;
	wire fragmenter_auto_out_d_valid;
	wire [2:0] fragmenter_auto_out_d_bits_opcode;
	wire [1:0] fragmenter_auto_out_d_bits_size;
	wire [7:0] fragmenter_auto_out_d_bits_source;
	wire [31:0] fragmenter_auto_out_d_bits_data;
	TLFragmenter_2 fragmenter(
		.clock(fragmenter_clock),
		.reset(fragmenter_reset),
		.auto_in_a_ready(fragmenter_auto_in_a_ready),
		.auto_in_a_valid(fragmenter_auto_in_a_valid),
		.auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
		.auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
		.auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
		.auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
		.auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
		.auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
		.auto_in_d_ready(fragmenter_auto_in_d_ready),
		.auto_in_d_valid(fragmenter_auto_in_d_valid),
		.auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
		.auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
		.auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
		.auto_out_a_ready(fragmenter_auto_out_a_ready),
		.auto_out_a_valid(fragmenter_auto_out_a_valid),
		.auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
		.auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
		.auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
		.auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
		.auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
		.auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
		.auto_out_d_ready(fragmenter_auto_out_d_ready),
		.auto_out_d_valid(fragmenter_auto_out_d_valid),
		.auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
		.auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
		.auto_out_d_bits_data(fragmenter_auto_out_d_bits_data)
	);
	assign auto_fragmenter_out_a_valid = fragmenter_auto_out_a_valid;
	assign auto_fragmenter_out_a_bits_opcode = fragmenter_auto_out_a_bits_opcode;
	assign auto_fragmenter_out_a_bits_param = fragmenter_auto_out_a_bits_param;
	assign auto_fragmenter_out_a_bits_size = fragmenter_auto_out_a_bits_size;
	assign auto_fragmenter_out_a_bits_source = fragmenter_auto_out_a_bits_source;
	assign auto_fragmenter_out_a_bits_address = fragmenter_auto_out_a_bits_address;
	assign auto_fragmenter_out_a_bits_mask = fragmenter_auto_out_a_bits_mask;
	assign auto_fragmenter_out_a_bits_data = fragmenter_auto_out_a_bits_data;
	assign auto_fragmenter_out_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt;
	assign auto_fragmenter_out_d_ready = fragmenter_auto_out_d_ready;
	assign auto_tl_in_a_ready = fragmenter_auto_in_a_ready;
	assign auto_tl_in_d_valid = fragmenter_auto_in_d_valid;
	assign auto_tl_in_d_bits_opcode = fragmenter_auto_in_d_bits_opcode;
	assign auto_tl_in_d_bits_size = fragmenter_auto_in_d_bits_size;
	assign auto_tl_in_d_bits_source = fragmenter_auto_in_d_bits_source;
	assign auto_tl_in_d_bits_data = fragmenter_auto_in_d_bits_data;
	assign fragmenter_clock = clock;
	assign fragmenter_reset = reset;
	assign fragmenter_auto_in_a_valid = auto_tl_in_a_valid;
	assign fragmenter_auto_in_a_bits_opcode = auto_tl_in_a_bits_opcode;
	assign fragmenter_auto_in_a_bits_param = auto_tl_in_a_bits_param;
	assign fragmenter_auto_in_a_bits_size = auto_tl_in_a_bits_size;
	assign fragmenter_auto_in_a_bits_source = auto_tl_in_a_bits_source;
	assign fragmenter_auto_in_a_bits_address = auto_tl_in_a_bits_address;
	assign fragmenter_auto_in_a_bits_mask = auto_tl_in_a_bits_mask;
	assign fragmenter_auto_in_a_bits_data = auto_tl_in_a_bits_data;
	assign fragmenter_auto_in_a_bits_corrupt = auto_tl_in_a_bits_corrupt;
	assign fragmenter_auto_in_d_ready = auto_tl_in_d_ready;
	assign fragmenter_auto_out_a_ready = auto_fragmenter_out_a_ready;
	assign fragmenter_auto_out_d_valid = auto_fragmenter_out_d_valid;
	assign fragmenter_auto_out_d_bits_opcode = auto_fragmenter_out_d_bits_opcode;
	assign fragmenter_auto_out_d_bits_size = auto_fragmenter_out_d_bits_size;
	assign fragmenter_auto_out_d_bits_source = auto_fragmenter_out_d_bits_source;
	assign fragmenter_auto_out_d_bits_data = auto_fragmenter_out_d_bits_data;
endmodule
module TLMonitor_24 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [25:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [25:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [25:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 26'h0000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [25:0] _T_56 = io_in_a_bits_address ^ 26'h2000000;
	wire [26:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [26:0] _T_59 = $signed(_T_57) & -27'sh0010000;
	wire _T_60 = $signed(_T_59) == 27'sh0000000;
	wire _T_92 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_96 = ~io_in_a_bits_mask;
	wire _T_97 = _T_96 == 4'h0;
	wire _T_101 = ~io_in_a_bits_corrupt;
	wire _T_105 = io_in_a_bits_opcode == 3'h7;
	wire _T_159 = io_in_a_bits_param != 3'h0;
	wire _T_172 = io_in_a_bits_opcode == 3'h4;
	wire _T_189 = io_in_a_bits_size <= 3'h6;
	wire _T_197 = _T_189 & _T_60;
	wire _T_208 = io_in_a_bits_param == 3'h0;
	wire _T_212 = io_in_a_bits_mask == mask;
	wire _T_220 = io_in_a_bits_opcode == 3'h0;
	wire _T_244 = source_ok & _T_197;
	wire _T_262 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_300 = ~mask;
	wire [3:0] _T_301 = io_in_a_bits_mask & _T_300;
	wire _T_302 = _T_301 == 4'h0;
	wire _T_306 = io_in_a_bits_opcode == 3'h2;
	wire _T_337 = io_in_a_bits_param <= 3'h4;
	wire _T_345 = io_in_a_bits_opcode == 3'h3;
	wire _T_376 = io_in_a_bits_param <= 3'h3;
	wire _T_384 = io_in_a_bits_opcode == 3'h5;
	wire _T_415 = io_in_a_bits_param <= 3'h1;
	wire _T_427 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_431 = io_in_d_bits_opcode == 3'h6;
	wire _T_435 = io_in_d_bits_size >= 3'h2;
	wire _T_451 = io_in_d_bits_opcode == 3'h4;
	wire _T_479 = io_in_d_bits_opcode == 3'h5;
	wire _T_508 = io_in_d_bits_opcode == 3'h0;
	wire _T_525 = io_in_d_bits_opcode == 3'h1;
	wire _T_543 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [25:0] address;
	wire _T_573 = io_in_a_valid & ~a_first;
	wire _T_574 = io_in_a_bits_opcode == opcode;
	wire _T_578 = io_in_a_bits_param == param;
	wire _T_582 = io_in_a_bits_size == size;
	wire _T_586 = io_in_a_bits_source == source;
	wire _T_590 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	wire _T_597 = io_in_d_valid & ~d_first;
	wire _T_598 = io_in_d_bits_opcode == opcode_1;
	wire _T_606 = io_in_d_bits_size == size_1;
	wire _T_610 = io_in_d_bits_source == source_1;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_624 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire _T_627 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_629 = inflight >> io_in_a_bits_source;
	wire _T_631 = ~_T_629[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_635 = io_in_d_valid & d_first_1;
	wire _T_637 = ~_T_431;
	wire _T_638 = (io_in_d_valid & d_first_1) & ~_T_431;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_637 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_637 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_624 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_648 = inflight >> io_in_d_bits_source;
	wire _T_650 = _T_648[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_655 = io_in_d_bits_opcode == _GEN_40;
	wire _T_656 = (io_in_d_bits_opcode == _GEN_32) | _T_655;
	wire _T_660 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_667 = io_in_d_bits_opcode == _GEN_56;
	wire _T_668 = (io_in_d_bits_opcode == _GEN_48) | _T_667;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_672 = _GEN_82 == a_size_lookup;
	wire _T_682 = (((_T_635 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_637;
	wire _T_684 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_693 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_719 = (io_in_d_valid & d_first_2) & _T_431;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_431 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_431 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_727 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_737 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_757 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Repeater_4 (
	clock,
	reset,
	io_repeat,
	io_full,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	input io_repeat;
	output wire io_full;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [25:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [25:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire io_deq_bits_corrupt;
	reg full;
	reg [2:0] saved_opcode;
	reg [2:0] saved_param;
	reg [2:0] saved_size;
	reg [2:0] saved_source;
	reg [25:0] saved_address;
	reg [3:0] saved_mask;
	reg saved_corrupt;
	wire _T = io_enq_ready & io_enq_valid;
	wire _GEN_0 = (_T & io_repeat) | full;
	wire _T_2 = io_deq_ready & io_deq_valid;
	assign io_full = full;
	assign io_enq_ready = io_deq_ready & ~full;
	assign io_deq_valid = io_enq_valid | full;
	assign io_deq_bits_opcode = (full ? saved_opcode : io_enq_bits_opcode);
	assign io_deq_bits_param = (full ? saved_param : io_enq_bits_param);
	assign io_deq_bits_size = (full ? saved_size : io_enq_bits_size);
	assign io_deq_bits_source = (full ? saved_source : io_enq_bits_source);
	assign io_deq_bits_address = (full ? saved_address : io_enq_bits_address);
	assign io_deq_bits_mask = (full ? saved_mask : io_enq_bits_mask);
	assign io_deq_bits_corrupt = (full ? saved_corrupt : io_enq_bits_corrupt);
	always @(posedge clock) begin
		if (reset)
			full <= 1'h0;
		else if (_T_2 & ~io_repeat)
			full <= 1'h0;
		else
			full <= _GEN_0;
		if (_T & io_repeat)
			saved_opcode <= io_enq_bits_opcode;
		if (_T & io_repeat)
			saved_param <= io_enq_bits_param;
		if (_T & io_repeat)
			saved_size <= io_enq_bits_size;
		if (_T & io_repeat)
			saved_source <= io_enq_bits_source;
		if (_T & io_repeat)
			saved_address <= io_enq_bits_address;
		if (_T & io_repeat)
			saved_mask <= io_enq_bits_mask;
		if (_T & io_repeat)
			saved_corrupt <= io_enq_bits_corrupt;
	end
endmodule
module TLFragmenter_3 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [25:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire [7:0] auto_out_a_bits_source;
	output wire [25:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_size;
	input [7:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [25:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire repeater_clock;
	wire repeater_reset;
	wire repeater_io_repeat;
	wire repeater_io_full;
	wire repeater_io_enq_ready;
	wire repeater_io_enq_valid;
	wire [2:0] repeater_io_enq_bits_opcode;
	wire [2:0] repeater_io_enq_bits_param;
	wire [2:0] repeater_io_enq_bits_size;
	wire [2:0] repeater_io_enq_bits_source;
	wire [25:0] repeater_io_enq_bits_address;
	wire [3:0] repeater_io_enq_bits_mask;
	wire repeater_io_enq_bits_corrupt;
	wire repeater_io_deq_ready;
	wire repeater_io_deq_valid;
	wire [2:0] repeater_io_deq_bits_opcode;
	wire [2:0] repeater_io_deq_bits_param;
	wire [2:0] repeater_io_deq_bits_size;
	wire [2:0] repeater_io_deq_bits_source;
	wire [25:0] repeater_io_deq_bits_address;
	wire [3:0] repeater_io_deq_bits_mask;
	wire repeater_io_deq_bits_corrupt;
	reg [3:0] acknum;
	reg [2:0] dOrig;
	reg dToggle;
	wire [3:0] dFragnum = auto_out_d_bits_source[3:0];
	wire dFirst = acknum == 4'h0;
	wire dLast = dFragnum == 4'h0;
	wire [3:0] _dsizeOH_T = 4'h1 << auto_out_d_bits_size;
	wire [2:0] dsizeOH = _dsizeOH_T[2:0];
	wire [4:0] _dsizeOH1_T_1 = 5'h03 << auto_out_d_bits_size;
	wire [1:0] dsizeOH1 = ~_dsizeOH1_T_1[1:0];
	wire dHasData = auto_out_d_bits_opcode[0];
	wire _T_5 = ~reset;
	wire ack_decrement = dHasData | dsizeOH[2];
	wire [5:0] _dFirst_size_T = {dFragnum, 2'h0};
	wire [5:0] _GEN_7 = {4'd0, dsizeOH1};
	wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7;
	wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0};
	wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h01;
	wire [6:0] _dFirst_size_T_4 = {1'h0, _dFirst_size_T_1};
	wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4;
	wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5;
	wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4];
	wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0];
	wire _dFirst_size_T_7 = |dFirst_size_hi;
	wire [3:0] _GEN_8 = {1'd0, dFirst_size_hi};
	wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo;
	wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2];
	wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0];
	wire _dFirst_size_T_9 = |dFirst_size_hi_1;
	wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1;
	wire [2:0] dFirst_size = {_dFirst_size_T_7, _dFirst_size_T_9, _dFirst_size_T_10[1]};
	wire drop = ~dHasData & ~dLast;
	wire bundleOut_0_d_ready = auto_in_d_ready | drop;
	wire _T_7 = bundleOut_0_d_ready & auto_out_d_valid;
	wire [3:0] _GEN_9 = {3'd0, ack_decrement};
	wire [3:0] _acknum_T_1 = acknum - _GEN_9;
	wire [2:0] aFrag = (repeater_io_deq_bits_size > 3'h2 ? 3'h2 : repeater_io_deq_bits_size);
	wire [12:0] _aOrigOH1_T_1 = 13'h003f << repeater_io_deq_bits_size;
	wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0];
	wire [8:0] _aFragOH1_T_1 = 9'h003 << aFrag;
	wire [1:0] aFragOH1 = ~_aFragOH1_T_1[1:0];
	wire aHasData = ~repeater_io_deq_bits_opcode[2];
	reg [3:0] gennum;
	wire aFirst = gennum == 4'h0;
	wire [3:0] _old_gennum1_T_2 = gennum - 4'h1;
	wire [3:0] old_gennum1 = (aFirst ? aOrigOH1[5:2] : _old_gennum1_T_2);
	wire [3:0] _new_gennum_T = ~old_gennum1;
	wire [3:0] new_gennum = ~_new_gennum_T;
	reg aToggle_r;
	wire _GEN_5 = (aFirst ? dToggle : aToggle_r);
	wire aToggle = ~_GEN_5;
	wire bundleOut_0_a_valid = repeater_io_deq_valid;
	wire _T_8 = auto_out_a_ready & bundleOut_0_a_valid;
	wire _repeater_io_repeat_T = ~aHasData;
	wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 2'h0};
	wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1;
	wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1;
	wire [5:0] _GEN_10 = {4'd0, aFragOH1};
	wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10;
	wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h03;
	wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4;
	wire [25:0] _GEN_11 = {20'd0, _bundleOut_0_a_bits_address_T_5};
	wire [3:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source, aToggle};
	wire _T_9 = ~repeater_io_full;
	TLMonitor_24 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	Repeater_4 repeater(
		.clock(repeater_clock),
		.reset(repeater_reset),
		.io_repeat(repeater_io_repeat),
		.io_full(repeater_io_full),
		.io_enq_ready(repeater_io_enq_ready),
		.io_enq_valid(repeater_io_enq_valid),
		.io_enq_bits_opcode(repeater_io_enq_bits_opcode),
		.io_enq_bits_param(repeater_io_enq_bits_param),
		.io_enq_bits_size(repeater_io_enq_bits_size),
		.io_enq_bits_source(repeater_io_enq_bits_source),
		.io_enq_bits_address(repeater_io_enq_bits_address),
		.io_enq_bits_mask(repeater_io_enq_bits_mask),
		.io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
		.io_deq_ready(repeater_io_deq_ready),
		.io_deq_valid(repeater_io_deq_valid),
		.io_deq_bits_opcode(repeater_io_deq_bits_opcode),
		.io_deq_bits_param(repeater_io_deq_bits_param),
		.io_deq_bits_size(repeater_io_deq_bits_size),
		.io_deq_bits_source(repeater_io_deq_bits_source),
		.io_deq_bits_address(repeater_io_deq_bits_address),
		.io_deq_bits_mask(repeater_io_deq_bits_mask),
		.io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = repeater_io_enq_ready;
	assign auto_in_d_valid = auto_out_d_valid & ~drop;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign auto_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_out_a_valid = repeater_io_deq_valid;
	assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode;
	assign auto_out_a_bits_param = repeater_io_deq_bits_param;
	assign auto_out_a_bits_size = aFrag[1:0];
	assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi, new_gennum};
	assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11;
	assign auto_out_a_bits_mask = (repeater_io_full ? 4'hf : auto_in_a_bits_mask);
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready | drop;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = repeater_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid & ~drop;
	assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_io_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign repeater_clock = clock;
	assign repeater_reset = reset;
	assign repeater_io_repeat = ~aHasData & (new_gennum != 4'h0);
	assign repeater_io_enq_valid = auto_in_a_valid;
	assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign repeater_io_enq_bits_param = auto_in_a_bits_param;
	assign repeater_io_enq_bits_size = auto_in_a_bits_size;
	assign repeater_io_enq_bits_source = auto_in_a_bits_source;
	assign repeater_io_enq_bits_address = auto_in_a_bits_address;
	assign repeater_io_enq_bits_mask = auto_in_a_bits_mask;
	assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign repeater_io_deq_ready = auto_out_a_ready;
	always @(posedge clock) begin
		if (reset)
			acknum <= 4'h0;
		else if (_T_7)
			if (dFirst)
				acknum <= dFragnum;
			else
				acknum <= _acknum_T_1;
		if (_T_7)
			if (dFirst)
				dOrig <= dFirst_size;
		if (reset)
			dToggle <= 1'h0;
		else if (_T_7)
			if (dFirst)
				dToggle <= auto_out_d_bits_source[4];
		if (reset)
			gennum <= 4'h0;
		else if (_T_8)
			gennum <= new_gennum;
		if (aFirst)
			aToggle_r <= dToggle;
	end
endmodule
module TLInterconnectCoupler_11 (
	clock,
	reset,
	auto_fragmenter_out_a_ready,
	auto_fragmenter_out_a_valid,
	auto_fragmenter_out_a_bits_opcode,
	auto_fragmenter_out_a_bits_param,
	auto_fragmenter_out_a_bits_size,
	auto_fragmenter_out_a_bits_source,
	auto_fragmenter_out_a_bits_address,
	auto_fragmenter_out_a_bits_mask,
	auto_fragmenter_out_a_bits_data,
	auto_fragmenter_out_a_bits_corrupt,
	auto_fragmenter_out_d_ready,
	auto_fragmenter_out_d_valid,
	auto_fragmenter_out_d_bits_opcode,
	auto_fragmenter_out_d_bits_size,
	auto_fragmenter_out_d_bits_source,
	auto_fragmenter_out_d_bits_data,
	auto_tl_in_a_ready,
	auto_tl_in_a_valid,
	auto_tl_in_a_bits_opcode,
	auto_tl_in_a_bits_param,
	auto_tl_in_a_bits_size,
	auto_tl_in_a_bits_source,
	auto_tl_in_a_bits_address,
	auto_tl_in_a_bits_mask,
	auto_tl_in_a_bits_data,
	auto_tl_in_a_bits_corrupt,
	auto_tl_in_d_ready,
	auto_tl_in_d_valid,
	auto_tl_in_d_bits_opcode,
	auto_tl_in_d_bits_size,
	auto_tl_in_d_bits_source,
	auto_tl_in_d_bits_data
);
	input clock;
	input reset;
	input auto_fragmenter_out_a_ready;
	output wire auto_fragmenter_out_a_valid;
	output wire [2:0] auto_fragmenter_out_a_bits_opcode;
	output wire [2:0] auto_fragmenter_out_a_bits_param;
	output wire [1:0] auto_fragmenter_out_a_bits_size;
	output wire [7:0] auto_fragmenter_out_a_bits_source;
	output wire [25:0] auto_fragmenter_out_a_bits_address;
	output wire [3:0] auto_fragmenter_out_a_bits_mask;
	output wire [31:0] auto_fragmenter_out_a_bits_data;
	output wire auto_fragmenter_out_a_bits_corrupt;
	output wire auto_fragmenter_out_d_ready;
	input auto_fragmenter_out_d_valid;
	input [2:0] auto_fragmenter_out_d_bits_opcode;
	input [1:0] auto_fragmenter_out_d_bits_size;
	input [7:0] auto_fragmenter_out_d_bits_source;
	input [31:0] auto_fragmenter_out_d_bits_data;
	output wire auto_tl_in_a_ready;
	input auto_tl_in_a_valid;
	input [2:0] auto_tl_in_a_bits_opcode;
	input [2:0] auto_tl_in_a_bits_param;
	input [2:0] auto_tl_in_a_bits_size;
	input [2:0] auto_tl_in_a_bits_source;
	input [25:0] auto_tl_in_a_bits_address;
	input [3:0] auto_tl_in_a_bits_mask;
	input [31:0] auto_tl_in_a_bits_data;
	input auto_tl_in_a_bits_corrupt;
	input auto_tl_in_d_ready;
	output wire auto_tl_in_d_valid;
	output wire [2:0] auto_tl_in_d_bits_opcode;
	output wire [2:0] auto_tl_in_d_bits_size;
	output wire [2:0] auto_tl_in_d_bits_source;
	output wire [31:0] auto_tl_in_d_bits_data;
	wire fragmenter_clock;
	wire fragmenter_reset;
	wire fragmenter_auto_in_a_ready;
	wire fragmenter_auto_in_a_valid;
	wire [2:0] fragmenter_auto_in_a_bits_opcode;
	wire [2:0] fragmenter_auto_in_a_bits_param;
	wire [2:0] fragmenter_auto_in_a_bits_size;
	wire [2:0] fragmenter_auto_in_a_bits_source;
	wire [25:0] fragmenter_auto_in_a_bits_address;
	wire [3:0] fragmenter_auto_in_a_bits_mask;
	wire [31:0] fragmenter_auto_in_a_bits_data;
	wire fragmenter_auto_in_a_bits_corrupt;
	wire fragmenter_auto_in_d_ready;
	wire fragmenter_auto_in_d_valid;
	wire [2:0] fragmenter_auto_in_d_bits_opcode;
	wire [2:0] fragmenter_auto_in_d_bits_size;
	wire [2:0] fragmenter_auto_in_d_bits_source;
	wire [31:0] fragmenter_auto_in_d_bits_data;
	wire fragmenter_auto_out_a_ready;
	wire fragmenter_auto_out_a_valid;
	wire [2:0] fragmenter_auto_out_a_bits_opcode;
	wire [2:0] fragmenter_auto_out_a_bits_param;
	wire [1:0] fragmenter_auto_out_a_bits_size;
	wire [7:0] fragmenter_auto_out_a_bits_source;
	wire [25:0] fragmenter_auto_out_a_bits_address;
	wire [3:0] fragmenter_auto_out_a_bits_mask;
	wire [31:0] fragmenter_auto_out_a_bits_data;
	wire fragmenter_auto_out_a_bits_corrupt;
	wire fragmenter_auto_out_d_ready;
	wire fragmenter_auto_out_d_valid;
	wire [2:0] fragmenter_auto_out_d_bits_opcode;
	wire [1:0] fragmenter_auto_out_d_bits_size;
	wire [7:0] fragmenter_auto_out_d_bits_source;
	wire [31:0] fragmenter_auto_out_d_bits_data;
	TLFragmenter_3 fragmenter(
		.clock(fragmenter_clock),
		.reset(fragmenter_reset),
		.auto_in_a_ready(fragmenter_auto_in_a_ready),
		.auto_in_a_valid(fragmenter_auto_in_a_valid),
		.auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
		.auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
		.auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
		.auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
		.auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
		.auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
		.auto_in_d_ready(fragmenter_auto_in_d_ready),
		.auto_in_d_valid(fragmenter_auto_in_d_valid),
		.auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
		.auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
		.auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
		.auto_out_a_ready(fragmenter_auto_out_a_ready),
		.auto_out_a_valid(fragmenter_auto_out_a_valid),
		.auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
		.auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
		.auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
		.auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
		.auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
		.auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
		.auto_out_d_ready(fragmenter_auto_out_d_ready),
		.auto_out_d_valid(fragmenter_auto_out_d_valid),
		.auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
		.auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
		.auto_out_d_bits_data(fragmenter_auto_out_d_bits_data)
	);
	assign auto_fragmenter_out_a_valid = fragmenter_auto_out_a_valid;
	assign auto_fragmenter_out_a_bits_opcode = fragmenter_auto_out_a_bits_opcode;
	assign auto_fragmenter_out_a_bits_param = fragmenter_auto_out_a_bits_param;
	assign auto_fragmenter_out_a_bits_size = fragmenter_auto_out_a_bits_size;
	assign auto_fragmenter_out_a_bits_source = fragmenter_auto_out_a_bits_source;
	assign auto_fragmenter_out_a_bits_address = fragmenter_auto_out_a_bits_address;
	assign auto_fragmenter_out_a_bits_mask = fragmenter_auto_out_a_bits_mask;
	assign auto_fragmenter_out_a_bits_data = fragmenter_auto_out_a_bits_data;
	assign auto_fragmenter_out_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt;
	assign auto_fragmenter_out_d_ready = fragmenter_auto_out_d_ready;
	assign auto_tl_in_a_ready = fragmenter_auto_in_a_ready;
	assign auto_tl_in_d_valid = fragmenter_auto_in_d_valid;
	assign auto_tl_in_d_bits_opcode = fragmenter_auto_in_d_bits_opcode;
	assign auto_tl_in_d_bits_size = fragmenter_auto_in_d_bits_size;
	assign auto_tl_in_d_bits_source = fragmenter_auto_in_d_bits_source;
	assign auto_tl_in_d_bits_data = fragmenter_auto_in_d_bits_data;
	assign fragmenter_clock = clock;
	assign fragmenter_reset = reset;
	assign fragmenter_auto_in_a_valid = auto_tl_in_a_valid;
	assign fragmenter_auto_in_a_bits_opcode = auto_tl_in_a_bits_opcode;
	assign fragmenter_auto_in_a_bits_param = auto_tl_in_a_bits_param;
	assign fragmenter_auto_in_a_bits_size = auto_tl_in_a_bits_size;
	assign fragmenter_auto_in_a_bits_source = auto_tl_in_a_bits_source;
	assign fragmenter_auto_in_a_bits_address = auto_tl_in_a_bits_address;
	assign fragmenter_auto_in_a_bits_mask = auto_tl_in_a_bits_mask;
	assign fragmenter_auto_in_a_bits_data = auto_tl_in_a_bits_data;
	assign fragmenter_auto_in_a_bits_corrupt = auto_tl_in_a_bits_corrupt;
	assign fragmenter_auto_in_d_ready = auto_tl_in_d_ready;
	assign fragmenter_auto_out_a_ready = auto_fragmenter_out_a_ready;
	assign fragmenter_auto_out_d_valid = auto_fragmenter_out_d_valid;
	assign fragmenter_auto_out_d_bits_opcode = auto_fragmenter_out_d_bits_opcode;
	assign fragmenter_auto_out_d_bits_size = auto_fragmenter_out_d_bits_size;
	assign fragmenter_auto_out_d_bits_source = auto_fragmenter_out_d_bits_source;
	assign fragmenter_auto_out_d_bits_data = auto_fragmenter_out_d_bits_data;
endmodule
module TLMonitor_25 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [11:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [11:0] _GEN_71 = {6'd0, is_aligned_mask};
	wire [11:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 12'h000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire [12:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [12:0] _T_59 = $signed(_T_7) & 13'sh1000;
	wire _T_60 = $signed(_T_59) == 13'sh0000;
	wire _T_92 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_96 = ~io_in_a_bits_mask;
	wire _T_97 = _T_96 == 4'h0;
	wire _T_101 = ~io_in_a_bits_corrupt;
	wire _T_105 = io_in_a_bits_opcode == 3'h7;
	wire _T_159 = io_in_a_bits_param != 3'h0;
	wire _T_172 = io_in_a_bits_opcode == 3'h4;
	wire _T_189 = io_in_a_bits_size <= 3'h6;
	wire _T_197 = _T_189 & _T_60;
	wire _T_208 = io_in_a_bits_param == 3'h0;
	wire _T_212 = io_in_a_bits_mask == mask;
	wire _T_220 = io_in_a_bits_opcode == 3'h0;
	wire _T_244 = source_ok & _T_197;
	wire _T_262 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_300 = ~mask;
	wire [3:0] _T_301 = io_in_a_bits_mask & _T_300;
	wire _T_302 = _T_301 == 4'h0;
	wire _T_306 = io_in_a_bits_opcode == 3'h2;
	wire _T_337 = io_in_a_bits_param <= 3'h4;
	wire _T_345 = io_in_a_bits_opcode == 3'h3;
	wire _T_376 = io_in_a_bits_param <= 3'h3;
	wire _T_384 = io_in_a_bits_opcode == 3'h5;
	wire _T_415 = io_in_a_bits_param <= 3'h1;
	wire _T_427 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_431 = io_in_d_bits_opcode == 3'h6;
	wire _T_435 = io_in_d_bits_size >= 3'h2;
	wire _T_451 = io_in_d_bits_opcode == 3'h4;
	wire _T_479 = io_in_d_bits_opcode == 3'h5;
	wire _T_508 = io_in_d_bits_opcode == 3'h0;
	wire _T_525 = io_in_d_bits_opcode == 3'h1;
	wire _T_543 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [11:0] address;
	wire _T_573 = io_in_a_valid & ~a_first;
	wire _T_574 = io_in_a_bits_opcode == opcode;
	wire _T_578 = io_in_a_bits_param == param;
	wire _T_582 = io_in_a_bits_size == size;
	wire _T_586 = io_in_a_bits_source == source;
	wire _T_590 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	wire _T_597 = io_in_d_valid & ~d_first;
	wire _T_598 = io_in_d_bits_opcode == opcode_1;
	wire _T_606 = io_in_d_bits_size == size_1;
	wire _T_610 = io_in_d_bits_source == source_1;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_624 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire _T_627 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_629 = inflight >> io_in_a_bits_source;
	wire _T_631 = ~_T_629[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_635 = io_in_d_valid & d_first_1;
	wire _T_637 = ~_T_431;
	wire _T_638 = (io_in_d_valid & d_first_1) & ~_T_431;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_637 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_637 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_624 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_648 = inflight >> io_in_d_bits_source;
	wire _T_650 = _T_648[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_655 = io_in_d_bits_opcode == _GEN_40;
	wire _T_656 = (io_in_d_bits_opcode == _GEN_32) | _T_655;
	wire _T_660 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_667 = io_in_d_bits_opcode == _GEN_56;
	wire _T_668 = (io_in_d_bits_opcode == _GEN_48) | _T_667;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_672 = _GEN_82 == a_size_lookup;
	wire _T_682 = (((_T_635 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_637;
	wire _T_684 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_693 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_719 = (io_in_d_valid & d_first_2) & _T_431;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_431 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_431 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_727 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_737 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_757 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Repeater_5 (
	clock,
	reset,
	io_repeat,
	io_full,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	input io_repeat;
	output wire io_full;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [11:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [11:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire io_deq_bits_corrupt;
	reg full;
	reg [2:0] saved_opcode;
	reg [2:0] saved_param;
	reg [2:0] saved_size;
	reg [2:0] saved_source;
	reg [11:0] saved_address;
	reg [3:0] saved_mask;
	reg saved_corrupt;
	wire _T = io_enq_ready & io_enq_valid;
	wire _GEN_0 = (_T & io_repeat) | full;
	wire _T_2 = io_deq_ready & io_deq_valid;
	assign io_full = full;
	assign io_enq_ready = io_deq_ready & ~full;
	assign io_deq_valid = io_enq_valid | full;
	assign io_deq_bits_opcode = (full ? saved_opcode : io_enq_bits_opcode);
	assign io_deq_bits_param = (full ? saved_param : io_enq_bits_param);
	assign io_deq_bits_size = (full ? saved_size : io_enq_bits_size);
	assign io_deq_bits_source = (full ? saved_source : io_enq_bits_source);
	assign io_deq_bits_address = (full ? saved_address : io_enq_bits_address);
	assign io_deq_bits_mask = (full ? saved_mask : io_enq_bits_mask);
	assign io_deq_bits_corrupt = (full ? saved_corrupt : io_enq_bits_corrupt);
	always @(posedge clock) begin
		if (reset)
			full <= 1'h0;
		else if (_T_2 & ~io_repeat)
			full <= 1'h0;
		else
			full <= _GEN_0;
		if (_T & io_repeat)
			saved_opcode <= io_enq_bits_opcode;
		if (_T & io_repeat)
			saved_param <= io_enq_bits_param;
		if (_T & io_repeat)
			saved_size <= io_enq_bits_size;
		if (_T & io_repeat)
			saved_source <= io_enq_bits_source;
		if (_T & io_repeat)
			saved_address <= io_enq_bits_address;
		if (_T & io_repeat)
			saved_mask <= io_enq_bits_mask;
		if (_T & io_repeat)
			saved_corrupt <= io_enq_bits_corrupt;
	end
endmodule
module TLFragmenter_4 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [11:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire [7:0] auto_out_a_bits_source;
	output wire [11:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_size;
	input [7:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [11:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire repeater_clock;
	wire repeater_reset;
	wire repeater_io_repeat;
	wire repeater_io_full;
	wire repeater_io_enq_ready;
	wire repeater_io_enq_valid;
	wire [2:0] repeater_io_enq_bits_opcode;
	wire [2:0] repeater_io_enq_bits_param;
	wire [2:0] repeater_io_enq_bits_size;
	wire [2:0] repeater_io_enq_bits_source;
	wire [11:0] repeater_io_enq_bits_address;
	wire [3:0] repeater_io_enq_bits_mask;
	wire repeater_io_enq_bits_corrupt;
	wire repeater_io_deq_ready;
	wire repeater_io_deq_valid;
	wire [2:0] repeater_io_deq_bits_opcode;
	wire [2:0] repeater_io_deq_bits_param;
	wire [2:0] repeater_io_deq_bits_size;
	wire [2:0] repeater_io_deq_bits_source;
	wire [11:0] repeater_io_deq_bits_address;
	wire [3:0] repeater_io_deq_bits_mask;
	wire repeater_io_deq_bits_corrupt;
	reg [3:0] acknum;
	reg [2:0] dOrig;
	reg dToggle;
	wire [3:0] dFragnum = auto_out_d_bits_source[3:0];
	wire dFirst = acknum == 4'h0;
	wire dLast = dFragnum == 4'h0;
	wire [3:0] _dsizeOH_T = 4'h1 << auto_out_d_bits_size;
	wire [2:0] dsizeOH = _dsizeOH_T[2:0];
	wire [4:0] _dsizeOH1_T_1 = 5'h03 << auto_out_d_bits_size;
	wire [1:0] dsizeOH1 = ~_dsizeOH1_T_1[1:0];
	wire dHasData = auto_out_d_bits_opcode[0];
	wire _T_5 = ~reset;
	wire ack_decrement = dHasData | dsizeOH[2];
	wire [5:0] _dFirst_size_T = {dFragnum, 2'h0};
	wire [5:0] _GEN_7 = {4'd0, dsizeOH1};
	wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7;
	wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0};
	wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h01;
	wire [6:0] _dFirst_size_T_4 = {1'h0, _dFirst_size_T_1};
	wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4;
	wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5;
	wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4];
	wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0];
	wire _dFirst_size_T_7 = |dFirst_size_hi;
	wire [3:0] _GEN_8 = {1'd0, dFirst_size_hi};
	wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo;
	wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2];
	wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0];
	wire _dFirst_size_T_9 = |dFirst_size_hi_1;
	wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1;
	wire [2:0] dFirst_size = {_dFirst_size_T_7, _dFirst_size_T_9, _dFirst_size_T_10[1]};
	wire drop = ~dHasData & ~dLast;
	wire bundleOut_0_d_ready = auto_in_d_ready | drop;
	wire _T_7 = bundleOut_0_d_ready & auto_out_d_valid;
	wire [3:0] _GEN_9 = {3'd0, ack_decrement};
	wire [3:0] _acknum_T_1 = acknum - _GEN_9;
	wire [2:0] aFrag = (repeater_io_deq_bits_size > 3'h2 ? 3'h2 : repeater_io_deq_bits_size);
	wire [12:0] _aOrigOH1_T_1 = 13'h003f << repeater_io_deq_bits_size;
	wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0];
	wire [8:0] _aFragOH1_T_1 = 9'h003 << aFrag;
	wire [1:0] aFragOH1 = ~_aFragOH1_T_1[1:0];
	wire aHasData = ~repeater_io_deq_bits_opcode[2];
	reg [3:0] gennum;
	wire aFirst = gennum == 4'h0;
	wire [3:0] _old_gennum1_T_2 = gennum - 4'h1;
	wire [3:0] old_gennum1 = (aFirst ? aOrigOH1[5:2] : _old_gennum1_T_2);
	wire [3:0] _new_gennum_T = ~old_gennum1;
	wire [3:0] new_gennum = ~_new_gennum_T;
	reg aToggle_r;
	wire _GEN_5 = (aFirst ? dToggle : aToggle_r);
	wire aToggle = ~_GEN_5;
	wire bundleOut_0_a_valid = repeater_io_deq_valid;
	wire _T_8 = auto_out_a_ready & bundleOut_0_a_valid;
	wire _repeater_io_repeat_T = ~aHasData;
	wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 2'h0};
	wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1;
	wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1;
	wire [5:0] _GEN_10 = {4'd0, aFragOH1};
	wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10;
	wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h03;
	wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4;
	wire [11:0] _GEN_11 = {6'd0, _bundleOut_0_a_bits_address_T_5};
	wire [3:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source, aToggle};
	wire _T_9 = ~repeater_io_full;
	TLMonitor_25 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	Repeater_5 repeater(
		.clock(repeater_clock),
		.reset(repeater_reset),
		.io_repeat(repeater_io_repeat),
		.io_full(repeater_io_full),
		.io_enq_ready(repeater_io_enq_ready),
		.io_enq_valid(repeater_io_enq_valid),
		.io_enq_bits_opcode(repeater_io_enq_bits_opcode),
		.io_enq_bits_param(repeater_io_enq_bits_param),
		.io_enq_bits_size(repeater_io_enq_bits_size),
		.io_enq_bits_source(repeater_io_enq_bits_source),
		.io_enq_bits_address(repeater_io_enq_bits_address),
		.io_enq_bits_mask(repeater_io_enq_bits_mask),
		.io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
		.io_deq_ready(repeater_io_deq_ready),
		.io_deq_valid(repeater_io_deq_valid),
		.io_deq_bits_opcode(repeater_io_deq_bits_opcode),
		.io_deq_bits_param(repeater_io_deq_bits_param),
		.io_deq_bits_size(repeater_io_deq_bits_size),
		.io_deq_bits_source(repeater_io_deq_bits_source),
		.io_deq_bits_address(repeater_io_deq_bits_address),
		.io_deq_bits_mask(repeater_io_deq_bits_mask),
		.io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = repeater_io_enq_ready;
	assign auto_in_d_valid = auto_out_d_valid & ~drop;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign auto_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_out_a_valid = repeater_io_deq_valid;
	assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode;
	assign auto_out_a_bits_param = repeater_io_deq_bits_param;
	assign auto_out_a_bits_size = aFrag[1:0];
	assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi, new_gennum};
	assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11;
	assign auto_out_a_bits_mask = (repeater_io_full ? 4'hf : auto_in_a_bits_mask);
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready | drop;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = repeater_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid & ~drop;
	assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_io_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign repeater_clock = clock;
	assign repeater_reset = reset;
	assign repeater_io_repeat = ~aHasData & (new_gennum != 4'h0);
	assign repeater_io_enq_valid = auto_in_a_valid;
	assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign repeater_io_enq_bits_param = auto_in_a_bits_param;
	assign repeater_io_enq_bits_size = auto_in_a_bits_size;
	assign repeater_io_enq_bits_source = auto_in_a_bits_source;
	assign repeater_io_enq_bits_address = auto_in_a_bits_address;
	assign repeater_io_enq_bits_mask = auto_in_a_bits_mask;
	assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign repeater_io_deq_ready = auto_out_a_ready;
	always @(posedge clock) begin
		if (reset)
			acknum <= 4'h0;
		else if (_T_7)
			if (dFirst)
				acknum <= dFragnum;
			else
				acknum <= _acknum_T_1;
		if (_T_7)
			if (dFirst)
				dOrig <= dFirst_size;
		if (reset)
			dToggle <= 1'h0;
		else if (_T_7)
			if (dFirst)
				dToggle <= auto_out_d_bits_source[4];
		if (reset)
			gennum <= 4'h0;
		else if (_T_8)
			gennum <= new_gennum;
		if (aFirst)
			aToggle_r <= dToggle;
	end
endmodule
module TLInterconnectCoupler_12 (
	clock,
	reset,
	auto_fragmenter_out_a_ready,
	auto_fragmenter_out_a_valid,
	auto_fragmenter_out_a_bits_opcode,
	auto_fragmenter_out_a_bits_param,
	auto_fragmenter_out_a_bits_size,
	auto_fragmenter_out_a_bits_source,
	auto_fragmenter_out_a_bits_address,
	auto_fragmenter_out_a_bits_mask,
	auto_fragmenter_out_a_bits_data,
	auto_fragmenter_out_a_bits_corrupt,
	auto_fragmenter_out_d_ready,
	auto_fragmenter_out_d_valid,
	auto_fragmenter_out_d_bits_opcode,
	auto_fragmenter_out_d_bits_size,
	auto_fragmenter_out_d_bits_source,
	auto_fragmenter_out_d_bits_data,
	auto_tl_in_a_ready,
	auto_tl_in_a_valid,
	auto_tl_in_a_bits_opcode,
	auto_tl_in_a_bits_param,
	auto_tl_in_a_bits_size,
	auto_tl_in_a_bits_source,
	auto_tl_in_a_bits_address,
	auto_tl_in_a_bits_mask,
	auto_tl_in_a_bits_data,
	auto_tl_in_a_bits_corrupt,
	auto_tl_in_d_ready,
	auto_tl_in_d_valid,
	auto_tl_in_d_bits_opcode,
	auto_tl_in_d_bits_size,
	auto_tl_in_d_bits_source,
	auto_tl_in_d_bits_data
);
	input clock;
	input reset;
	input auto_fragmenter_out_a_ready;
	output wire auto_fragmenter_out_a_valid;
	output wire [2:0] auto_fragmenter_out_a_bits_opcode;
	output wire [2:0] auto_fragmenter_out_a_bits_param;
	output wire [1:0] auto_fragmenter_out_a_bits_size;
	output wire [7:0] auto_fragmenter_out_a_bits_source;
	output wire [11:0] auto_fragmenter_out_a_bits_address;
	output wire [3:0] auto_fragmenter_out_a_bits_mask;
	output wire [31:0] auto_fragmenter_out_a_bits_data;
	output wire auto_fragmenter_out_a_bits_corrupt;
	output wire auto_fragmenter_out_d_ready;
	input auto_fragmenter_out_d_valid;
	input [2:0] auto_fragmenter_out_d_bits_opcode;
	input [1:0] auto_fragmenter_out_d_bits_size;
	input [7:0] auto_fragmenter_out_d_bits_source;
	input [31:0] auto_fragmenter_out_d_bits_data;
	output wire auto_tl_in_a_ready;
	input auto_tl_in_a_valid;
	input [2:0] auto_tl_in_a_bits_opcode;
	input [2:0] auto_tl_in_a_bits_param;
	input [2:0] auto_tl_in_a_bits_size;
	input [2:0] auto_tl_in_a_bits_source;
	input [11:0] auto_tl_in_a_bits_address;
	input [3:0] auto_tl_in_a_bits_mask;
	input [31:0] auto_tl_in_a_bits_data;
	input auto_tl_in_a_bits_corrupt;
	input auto_tl_in_d_ready;
	output wire auto_tl_in_d_valid;
	output wire [2:0] auto_tl_in_d_bits_opcode;
	output wire [2:0] auto_tl_in_d_bits_size;
	output wire [2:0] auto_tl_in_d_bits_source;
	output wire [31:0] auto_tl_in_d_bits_data;
	wire fragmenter_clock;
	wire fragmenter_reset;
	wire fragmenter_auto_in_a_ready;
	wire fragmenter_auto_in_a_valid;
	wire [2:0] fragmenter_auto_in_a_bits_opcode;
	wire [2:0] fragmenter_auto_in_a_bits_param;
	wire [2:0] fragmenter_auto_in_a_bits_size;
	wire [2:0] fragmenter_auto_in_a_bits_source;
	wire [11:0] fragmenter_auto_in_a_bits_address;
	wire [3:0] fragmenter_auto_in_a_bits_mask;
	wire [31:0] fragmenter_auto_in_a_bits_data;
	wire fragmenter_auto_in_a_bits_corrupt;
	wire fragmenter_auto_in_d_ready;
	wire fragmenter_auto_in_d_valid;
	wire [2:0] fragmenter_auto_in_d_bits_opcode;
	wire [2:0] fragmenter_auto_in_d_bits_size;
	wire [2:0] fragmenter_auto_in_d_bits_source;
	wire [31:0] fragmenter_auto_in_d_bits_data;
	wire fragmenter_auto_out_a_ready;
	wire fragmenter_auto_out_a_valid;
	wire [2:0] fragmenter_auto_out_a_bits_opcode;
	wire [2:0] fragmenter_auto_out_a_bits_param;
	wire [1:0] fragmenter_auto_out_a_bits_size;
	wire [7:0] fragmenter_auto_out_a_bits_source;
	wire [11:0] fragmenter_auto_out_a_bits_address;
	wire [3:0] fragmenter_auto_out_a_bits_mask;
	wire [31:0] fragmenter_auto_out_a_bits_data;
	wire fragmenter_auto_out_a_bits_corrupt;
	wire fragmenter_auto_out_d_ready;
	wire fragmenter_auto_out_d_valid;
	wire [2:0] fragmenter_auto_out_d_bits_opcode;
	wire [1:0] fragmenter_auto_out_d_bits_size;
	wire [7:0] fragmenter_auto_out_d_bits_source;
	wire [31:0] fragmenter_auto_out_d_bits_data;
	TLFragmenter_4 fragmenter(
		.clock(fragmenter_clock),
		.reset(fragmenter_reset),
		.auto_in_a_ready(fragmenter_auto_in_a_ready),
		.auto_in_a_valid(fragmenter_auto_in_a_valid),
		.auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
		.auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
		.auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
		.auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
		.auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
		.auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
		.auto_in_d_ready(fragmenter_auto_in_d_ready),
		.auto_in_d_valid(fragmenter_auto_in_d_valid),
		.auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
		.auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
		.auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
		.auto_out_a_ready(fragmenter_auto_out_a_ready),
		.auto_out_a_valid(fragmenter_auto_out_a_valid),
		.auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
		.auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
		.auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
		.auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
		.auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
		.auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
		.auto_out_d_ready(fragmenter_auto_out_d_ready),
		.auto_out_d_valid(fragmenter_auto_out_d_valid),
		.auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
		.auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
		.auto_out_d_bits_data(fragmenter_auto_out_d_bits_data)
	);
	assign auto_fragmenter_out_a_valid = fragmenter_auto_out_a_valid;
	assign auto_fragmenter_out_a_bits_opcode = fragmenter_auto_out_a_bits_opcode;
	assign auto_fragmenter_out_a_bits_param = fragmenter_auto_out_a_bits_param;
	assign auto_fragmenter_out_a_bits_size = fragmenter_auto_out_a_bits_size;
	assign auto_fragmenter_out_a_bits_source = fragmenter_auto_out_a_bits_source;
	assign auto_fragmenter_out_a_bits_address = fragmenter_auto_out_a_bits_address;
	assign auto_fragmenter_out_a_bits_mask = fragmenter_auto_out_a_bits_mask;
	assign auto_fragmenter_out_a_bits_data = fragmenter_auto_out_a_bits_data;
	assign auto_fragmenter_out_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt;
	assign auto_fragmenter_out_d_ready = fragmenter_auto_out_d_ready;
	assign auto_tl_in_a_ready = fragmenter_auto_in_a_ready;
	assign auto_tl_in_d_valid = fragmenter_auto_in_d_valid;
	assign auto_tl_in_d_bits_opcode = fragmenter_auto_in_d_bits_opcode;
	assign auto_tl_in_d_bits_size = fragmenter_auto_in_d_bits_size;
	assign auto_tl_in_d_bits_source = fragmenter_auto_in_d_bits_source;
	assign auto_tl_in_d_bits_data = fragmenter_auto_in_d_bits_data;
	assign fragmenter_clock = clock;
	assign fragmenter_reset = reset;
	assign fragmenter_auto_in_a_valid = auto_tl_in_a_valid;
	assign fragmenter_auto_in_a_bits_opcode = auto_tl_in_a_bits_opcode;
	assign fragmenter_auto_in_a_bits_param = auto_tl_in_a_bits_param;
	assign fragmenter_auto_in_a_bits_size = auto_tl_in_a_bits_size;
	assign fragmenter_auto_in_a_bits_source = auto_tl_in_a_bits_source;
	assign fragmenter_auto_in_a_bits_address = auto_tl_in_a_bits_address;
	assign fragmenter_auto_in_a_bits_mask = auto_tl_in_a_bits_mask;
	assign fragmenter_auto_in_a_bits_data = auto_tl_in_a_bits_data;
	assign fragmenter_auto_in_a_bits_corrupt = auto_tl_in_a_bits_corrupt;
	assign fragmenter_auto_in_d_ready = auto_tl_in_d_ready;
	assign fragmenter_auto_out_a_ready = auto_fragmenter_out_a_ready;
	assign fragmenter_auto_out_d_valid = auto_fragmenter_out_d_valid;
	assign fragmenter_auto_out_d_bits_opcode = auto_fragmenter_out_d_bits_opcode;
	assign fragmenter_auto_out_d_bits_size = auto_fragmenter_out_d_bits_size;
	assign fragmenter_auto_out_d_bits_source = auto_fragmenter_out_d_bits_source;
	assign fragmenter_auto_out_d_bits_data = auto_fragmenter_out_d_bits_data;
endmodule
module TLWidthWidget_6 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module TLInterconnectCoupler_13 (
	auto_tl_slave_clock_xing_out_a_ready,
	auto_tl_slave_clock_xing_out_a_valid,
	auto_tl_slave_clock_xing_out_a_bits_opcode,
	auto_tl_slave_clock_xing_out_a_bits_param,
	auto_tl_slave_clock_xing_out_a_bits_size,
	auto_tl_slave_clock_xing_out_a_bits_source,
	auto_tl_slave_clock_xing_out_a_bits_address,
	auto_tl_slave_clock_xing_out_a_bits_mask,
	auto_tl_slave_clock_xing_out_a_bits_data,
	auto_tl_slave_clock_xing_out_d_ready,
	auto_tl_slave_clock_xing_out_d_valid,
	auto_tl_slave_clock_xing_out_d_bits_opcode,
	auto_tl_slave_clock_xing_out_d_bits_param,
	auto_tl_slave_clock_xing_out_d_bits_size,
	auto_tl_slave_clock_xing_out_d_bits_source,
	auto_tl_slave_clock_xing_out_d_bits_sink,
	auto_tl_slave_clock_xing_out_d_bits_denied,
	auto_tl_slave_clock_xing_out_d_bits_data,
	auto_tl_slave_clock_xing_out_d_bits_corrupt,
	auto_tl_in_a_ready,
	auto_tl_in_a_valid,
	auto_tl_in_a_bits_opcode,
	auto_tl_in_a_bits_param,
	auto_tl_in_a_bits_size,
	auto_tl_in_a_bits_source,
	auto_tl_in_a_bits_address,
	auto_tl_in_a_bits_mask,
	auto_tl_in_a_bits_data,
	auto_tl_in_d_ready,
	auto_tl_in_d_valid,
	auto_tl_in_d_bits_opcode,
	auto_tl_in_d_bits_param,
	auto_tl_in_d_bits_size,
	auto_tl_in_d_bits_source,
	auto_tl_in_d_bits_sink,
	auto_tl_in_d_bits_denied,
	auto_tl_in_d_bits_data,
	auto_tl_in_d_bits_corrupt
);
	input auto_tl_slave_clock_xing_out_a_ready;
	output wire auto_tl_slave_clock_xing_out_a_valid;
	output wire [2:0] auto_tl_slave_clock_xing_out_a_bits_opcode;
	output wire [2:0] auto_tl_slave_clock_xing_out_a_bits_param;
	output wire [2:0] auto_tl_slave_clock_xing_out_a_bits_size;
	output wire [2:0] auto_tl_slave_clock_xing_out_a_bits_source;
	output wire [31:0] auto_tl_slave_clock_xing_out_a_bits_address;
	output wire [3:0] auto_tl_slave_clock_xing_out_a_bits_mask;
	output wire [31:0] auto_tl_slave_clock_xing_out_a_bits_data;
	output wire auto_tl_slave_clock_xing_out_d_ready;
	input auto_tl_slave_clock_xing_out_d_valid;
	input [2:0] auto_tl_slave_clock_xing_out_d_bits_opcode;
	input [1:0] auto_tl_slave_clock_xing_out_d_bits_param;
	input [2:0] auto_tl_slave_clock_xing_out_d_bits_size;
	input [2:0] auto_tl_slave_clock_xing_out_d_bits_source;
	input auto_tl_slave_clock_xing_out_d_bits_sink;
	input auto_tl_slave_clock_xing_out_d_bits_denied;
	input [31:0] auto_tl_slave_clock_xing_out_d_bits_data;
	input auto_tl_slave_clock_xing_out_d_bits_corrupt;
	output wire auto_tl_in_a_ready;
	input auto_tl_in_a_valid;
	input [2:0] auto_tl_in_a_bits_opcode;
	input [2:0] auto_tl_in_a_bits_param;
	input [2:0] auto_tl_in_a_bits_size;
	input [2:0] auto_tl_in_a_bits_source;
	input [31:0] auto_tl_in_a_bits_address;
	input [3:0] auto_tl_in_a_bits_mask;
	input [31:0] auto_tl_in_a_bits_data;
	input auto_tl_in_d_ready;
	output wire auto_tl_in_d_valid;
	output wire [2:0] auto_tl_in_d_bits_opcode;
	output wire [1:0] auto_tl_in_d_bits_param;
	output wire [2:0] auto_tl_in_d_bits_size;
	output wire [2:0] auto_tl_in_d_bits_source;
	output wire auto_tl_in_d_bits_sink;
	output wire auto_tl_in_d_bits_denied;
	output wire [31:0] auto_tl_in_d_bits_data;
	output wire auto_tl_in_d_bits_corrupt;
	wire widget_auto_in_a_ready;
	wire widget_auto_in_a_valid;
	wire [2:0] widget_auto_in_a_bits_opcode;
	wire [2:0] widget_auto_in_a_bits_param;
	wire [2:0] widget_auto_in_a_bits_size;
	wire [2:0] widget_auto_in_a_bits_source;
	wire [31:0] widget_auto_in_a_bits_address;
	wire [3:0] widget_auto_in_a_bits_mask;
	wire [31:0] widget_auto_in_a_bits_data;
	wire widget_auto_in_d_ready;
	wire widget_auto_in_d_valid;
	wire [2:0] widget_auto_in_d_bits_opcode;
	wire [1:0] widget_auto_in_d_bits_param;
	wire [2:0] widget_auto_in_d_bits_size;
	wire [2:0] widget_auto_in_d_bits_source;
	wire widget_auto_in_d_bits_sink;
	wire widget_auto_in_d_bits_denied;
	wire [31:0] widget_auto_in_d_bits_data;
	wire widget_auto_in_d_bits_corrupt;
	wire widget_auto_out_a_ready;
	wire widget_auto_out_a_valid;
	wire [2:0] widget_auto_out_a_bits_opcode;
	wire [2:0] widget_auto_out_a_bits_param;
	wire [2:0] widget_auto_out_a_bits_size;
	wire [2:0] widget_auto_out_a_bits_source;
	wire [31:0] widget_auto_out_a_bits_address;
	wire [3:0] widget_auto_out_a_bits_mask;
	wire [31:0] widget_auto_out_a_bits_data;
	wire widget_auto_out_d_ready;
	wire widget_auto_out_d_valid;
	wire [2:0] widget_auto_out_d_bits_opcode;
	wire [1:0] widget_auto_out_d_bits_param;
	wire [2:0] widget_auto_out_d_bits_size;
	wire [2:0] widget_auto_out_d_bits_source;
	wire widget_auto_out_d_bits_sink;
	wire widget_auto_out_d_bits_denied;
	wire [31:0] widget_auto_out_d_bits_data;
	wire widget_auto_out_d_bits_corrupt;
	TLWidthWidget_6 widget(
		.auto_in_a_ready(widget_auto_in_a_ready),
		.auto_in_a_valid(widget_auto_in_a_valid),
		.auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(widget_auto_in_a_bits_param),
		.auto_in_a_bits_size(widget_auto_in_a_bits_size),
		.auto_in_a_bits_source(widget_auto_in_a_bits_source),
		.auto_in_a_bits_address(widget_auto_in_a_bits_address),
		.auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
		.auto_in_a_bits_data(widget_auto_in_a_bits_data),
		.auto_in_d_ready(widget_auto_in_d_ready),
		.auto_in_d_valid(widget_auto_in_d_valid),
		.auto_in_d_bits_opcode(widget_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(widget_auto_in_d_bits_param),
		.auto_in_d_bits_size(widget_auto_in_d_bits_size),
		.auto_in_d_bits_source(widget_auto_in_d_bits_source),
		.auto_in_d_bits_sink(widget_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(widget_auto_in_d_bits_denied),
		.auto_in_d_bits_data(widget_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(widget_auto_in_d_bits_corrupt),
		.auto_out_a_ready(widget_auto_out_a_ready),
		.auto_out_a_valid(widget_auto_out_a_valid),
		.auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(widget_auto_out_a_bits_param),
		.auto_out_a_bits_size(widget_auto_out_a_bits_size),
		.auto_out_a_bits_source(widget_auto_out_a_bits_source),
		.auto_out_a_bits_address(widget_auto_out_a_bits_address),
		.auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
		.auto_out_a_bits_data(widget_auto_out_a_bits_data),
		.auto_out_d_ready(widget_auto_out_d_ready),
		.auto_out_d_valid(widget_auto_out_d_valid),
		.auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(widget_auto_out_d_bits_param),
		.auto_out_d_bits_size(widget_auto_out_d_bits_size),
		.auto_out_d_bits_source(widget_auto_out_d_bits_source),
		.auto_out_d_bits_sink(widget_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(widget_auto_out_d_bits_denied),
		.auto_out_d_bits_data(widget_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(widget_auto_out_d_bits_corrupt)
	);
	assign auto_tl_slave_clock_xing_out_a_valid = widget_auto_out_a_valid;
	assign auto_tl_slave_clock_xing_out_a_bits_opcode = widget_auto_out_a_bits_opcode;
	assign auto_tl_slave_clock_xing_out_a_bits_param = widget_auto_out_a_bits_param;
	assign auto_tl_slave_clock_xing_out_a_bits_size = widget_auto_out_a_bits_size;
	assign auto_tl_slave_clock_xing_out_a_bits_source = widget_auto_out_a_bits_source;
	assign auto_tl_slave_clock_xing_out_a_bits_address = widget_auto_out_a_bits_address;
	assign auto_tl_slave_clock_xing_out_a_bits_mask = widget_auto_out_a_bits_mask;
	assign auto_tl_slave_clock_xing_out_a_bits_data = widget_auto_out_a_bits_data;
	assign auto_tl_slave_clock_xing_out_d_ready = widget_auto_out_d_ready;
	assign auto_tl_in_a_ready = widget_auto_in_a_ready;
	assign auto_tl_in_d_valid = widget_auto_in_d_valid;
	assign auto_tl_in_d_bits_opcode = widget_auto_in_d_bits_opcode;
	assign auto_tl_in_d_bits_param = widget_auto_in_d_bits_param;
	assign auto_tl_in_d_bits_size = widget_auto_in_d_bits_size;
	assign auto_tl_in_d_bits_source = widget_auto_in_d_bits_source;
	assign auto_tl_in_d_bits_sink = widget_auto_in_d_bits_sink;
	assign auto_tl_in_d_bits_denied = widget_auto_in_d_bits_denied;
	assign auto_tl_in_d_bits_data = widget_auto_in_d_bits_data;
	assign auto_tl_in_d_bits_corrupt = widget_auto_in_d_bits_corrupt;
	assign widget_auto_in_a_valid = auto_tl_in_a_valid;
	assign widget_auto_in_a_bits_opcode = auto_tl_in_a_bits_opcode;
	assign widget_auto_in_a_bits_param = auto_tl_in_a_bits_param;
	assign widget_auto_in_a_bits_size = auto_tl_in_a_bits_size;
	assign widget_auto_in_a_bits_source = auto_tl_in_a_bits_source;
	assign widget_auto_in_a_bits_address = auto_tl_in_a_bits_address;
	assign widget_auto_in_a_bits_mask = auto_tl_in_a_bits_mask;
	assign widget_auto_in_a_bits_data = auto_tl_in_a_bits_data;
	assign widget_auto_in_d_ready = auto_tl_in_d_ready;
	assign widget_auto_out_a_ready = auto_tl_slave_clock_xing_out_a_ready;
	assign widget_auto_out_d_valid = auto_tl_slave_clock_xing_out_d_valid;
	assign widget_auto_out_d_bits_opcode = auto_tl_slave_clock_xing_out_d_bits_opcode;
	assign widget_auto_out_d_bits_param = auto_tl_slave_clock_xing_out_d_bits_param;
	assign widget_auto_out_d_bits_size = auto_tl_slave_clock_xing_out_d_bits_size;
	assign widget_auto_out_d_bits_source = auto_tl_slave_clock_xing_out_d_bits_source;
	assign widget_auto_out_d_bits_sink = auto_tl_slave_clock_xing_out_d_bits_sink;
	assign widget_auto_out_d_bits_denied = auto_tl_slave_clock_xing_out_d_bits_denied;
	assign widget_auto_out_d_bits_data = auto_tl_slave_clock_xing_out_d_bits_data;
	assign widget_auto_out_d_bits_corrupt = auto_tl_slave_clock_xing_out_d_bits_corrupt;
endmodule
module TLMonitor_26 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [16:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [16:0] _GEN_71 = {11'd0, is_aligned_mask};
	wire [16:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 17'h00000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [16:0] _T_56 = io_in_a_bits_address ^ 17'h10000;
	wire [17:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [17:0] _T_59 = $signed(_T_57) & -18'sh10000;
	wire _T_60 = $signed(_T_59) == 18'sh00000;
	wire _T_92 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_96 = ~io_in_a_bits_mask;
	wire _T_97 = _T_96 == 4'h0;
	wire _T_101 = ~io_in_a_bits_corrupt;
	wire _T_105 = io_in_a_bits_opcode == 3'h7;
	wire _T_159 = io_in_a_bits_param != 3'h0;
	wire _T_172 = io_in_a_bits_opcode == 3'h4;
	wire _T_189 = io_in_a_bits_size <= 3'h6;
	wire _T_197 = _T_189 & _T_60;
	wire _T_208 = io_in_a_bits_param == 3'h0;
	wire _T_212 = io_in_a_bits_mask == mask;
	wire _T_220 = io_in_a_bits_opcode == 3'h0;
	wire _T_259 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_294 = ~mask;
	wire [3:0] _T_295 = io_in_a_bits_mask & _T_294;
	wire _T_296 = _T_295 == 4'h0;
	wire _T_300 = io_in_a_bits_opcode == 3'h2;
	wire _T_331 = io_in_a_bits_param <= 3'h4;
	wire _T_339 = io_in_a_bits_opcode == 3'h3;
	wire _T_370 = io_in_a_bits_param <= 3'h3;
	wire _T_378 = io_in_a_bits_opcode == 3'h5;
	wire _T_409 = io_in_a_bits_param <= 3'h1;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [16:0] address;
	wire _T_567 = io_in_a_valid & ~a_first;
	wire _T_568 = io_in_a_bits_opcode == opcode;
	wire _T_572 = io_in_a_bits_param == param;
	wire _T_576 = io_in_a_bits_size == size;
	wire _T_580 = io_in_a_bits_source == source;
	wire _T_584 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] size_1;
	reg [2:0] source_1;
	wire _T_591 = io_in_d_valid & ~d_first;
	wire _T_600 = io_in_d_bits_size == size_1;
	wire _T_604 = io_in_d_bits_source == source_1;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_618 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire _T_621 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (a_first_done & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_623 = inflight >> io_in_a_bits_source;
	wire _T_625 = ~_T_623[0];
	wire [7:0] _GEN_16 = (a_first_done & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_629 = io_in_d_valid & d_first_1;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = (_d_first_T & d_first_1 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = (_d_first_T & d_first_1 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_618 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_642 = inflight >> io_in_d_bits_source;
	wire _T_644 = _T_642[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_649 = 3'h1 == _GEN_40;
	wire _T_650 = (3'h1 == _GEN_32) | _T_649;
	wire _T_654 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_661 = 3'h1 == _GEN_56;
	wire _T_662 = (3'h1 == _GEN_48) | _T_661;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_666 = _GEN_82 == a_size_lookup;
	wire _T_674 = ((_T_629 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2;
	wire _T_678 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_687 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 4'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			param <= io_in_a_bits_param;
		if (a_first_done & a_first)
			size <= io_in_a_bits_size;
		if (a_first_done & a_first)
			source <= io_in_a_bits_source;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first)
				d_first_counter <= d_first_beats1_decode;
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 4'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1)
				d_first_counter_1 <= d_first_beats1_decode;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
	end
endmodule
module Repeater_6 (
	clock,
	reset,
	io_repeat,
	io_full,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	input io_repeat;
	output wire io_full;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [16:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [16:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire io_deq_bits_corrupt;
	reg full;
	reg [2:0] saved_opcode;
	reg [2:0] saved_param;
	reg [2:0] saved_size;
	reg [2:0] saved_source;
	reg [16:0] saved_address;
	reg [3:0] saved_mask;
	reg saved_corrupt;
	wire _T = io_enq_ready & io_enq_valid;
	wire _GEN_0 = (_T & io_repeat) | full;
	wire _T_2 = io_deq_ready & io_deq_valid;
	assign io_full = full;
	assign io_enq_ready = io_deq_ready & ~full;
	assign io_deq_valid = io_enq_valid | full;
	assign io_deq_bits_opcode = (full ? saved_opcode : io_enq_bits_opcode);
	assign io_deq_bits_param = (full ? saved_param : io_enq_bits_param);
	assign io_deq_bits_size = (full ? saved_size : io_enq_bits_size);
	assign io_deq_bits_source = (full ? saved_source : io_enq_bits_source);
	assign io_deq_bits_address = (full ? saved_address : io_enq_bits_address);
	assign io_deq_bits_mask = (full ? saved_mask : io_enq_bits_mask);
	assign io_deq_bits_corrupt = (full ? saved_corrupt : io_enq_bits_corrupt);
	always @(posedge clock) begin
		if (reset)
			full <= 1'h0;
		else if (_T_2 & ~io_repeat)
			full <= 1'h0;
		else
			full <= _GEN_0;
		if (_T & io_repeat)
			saved_opcode <= io_enq_bits_opcode;
		if (_T & io_repeat)
			saved_param <= io_enq_bits_param;
		if (_T & io_repeat)
			saved_size <= io_enq_bits_size;
		if (_T & io_repeat)
			saved_source <= io_enq_bits_source;
		if (_T & io_repeat)
			saved_address <= io_enq_bits_address;
		if (_T & io_repeat)
			saved_mask <= io_enq_bits_mask;
		if (_T & io_repeat)
			saved_corrupt <= io_enq_bits_corrupt;
	end
endmodule
module TLFragmenter_5 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [16:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire [7:0] auto_out_a_bits_source;
	output wire [16:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [1:0] auto_out_d_bits_size;
	input [7:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [16:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire repeater_clock;
	wire repeater_reset;
	wire repeater_io_repeat;
	wire repeater_io_full;
	wire repeater_io_enq_ready;
	wire repeater_io_enq_valid;
	wire [2:0] repeater_io_enq_bits_opcode;
	wire [2:0] repeater_io_enq_bits_param;
	wire [2:0] repeater_io_enq_bits_size;
	wire [2:0] repeater_io_enq_bits_source;
	wire [16:0] repeater_io_enq_bits_address;
	wire [3:0] repeater_io_enq_bits_mask;
	wire repeater_io_enq_bits_corrupt;
	wire repeater_io_deq_ready;
	wire repeater_io_deq_valid;
	wire [2:0] repeater_io_deq_bits_opcode;
	wire [2:0] repeater_io_deq_bits_param;
	wire [2:0] repeater_io_deq_bits_size;
	wire [2:0] repeater_io_deq_bits_source;
	wire [16:0] repeater_io_deq_bits_address;
	wire [3:0] repeater_io_deq_bits_mask;
	wire repeater_io_deq_bits_corrupt;
	reg [3:0] acknum;
	reg [2:0] dOrig;
	reg dToggle;
	wire [3:0] dFragnum = auto_out_d_bits_source[3:0];
	wire dFirst = acknum == 4'h0;
	wire [4:0] _dsizeOH1_T_1 = 5'h03 << auto_out_d_bits_size;
	wire [1:0] dsizeOH1 = ~_dsizeOH1_T_1[1:0];
	wire _T_5 = ~reset;
	wire [5:0] _dFirst_size_T = {dFragnum, 2'h0};
	wire [5:0] _GEN_7 = {4'd0, dsizeOH1};
	wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7;
	wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0};
	wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h01;
	wire [6:0] _dFirst_size_T_4 = {1'h0, _dFirst_size_T_1};
	wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4;
	wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5;
	wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4];
	wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0];
	wire _dFirst_size_T_7 = |dFirst_size_hi;
	wire [3:0] _GEN_8 = {1'd0, dFirst_size_hi};
	wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo;
	wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2];
	wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0];
	wire _dFirst_size_T_9 = |dFirst_size_hi_1;
	wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1;
	wire [2:0] dFirst_size = {_dFirst_size_T_7, _dFirst_size_T_9, _dFirst_size_T_10[1]};
	wire _T_7 = auto_in_d_ready & auto_out_d_valid;
	wire [3:0] _acknum_T_1 = acknum - 4'h1;
	wire [2:0] aFrag = (repeater_io_deq_bits_size > 3'h2 ? 3'h2 : repeater_io_deq_bits_size);
	wire [12:0] _aOrigOH1_T_1 = 13'h003f << repeater_io_deq_bits_size;
	wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0];
	wire [8:0] _aFragOH1_T_1 = 9'h003 << aFrag;
	wire [1:0] aFragOH1 = ~_aFragOH1_T_1[1:0];
	reg [3:0] gennum;
	wire aFirst = gennum == 4'h0;
	wire [3:0] _old_gennum1_T_2 = gennum - 4'h1;
	wire [3:0] old_gennum1 = (aFirst ? aOrigOH1[5:2] : _old_gennum1_T_2);
	wire [3:0] _new_gennum_T = ~old_gennum1;
	wire [3:0] new_gennum = ~_new_gennum_T;
	reg aToggle_r;
	wire _GEN_5 = (aFirst ? dToggle : aToggle_r);
	wire aToggle = ~_GEN_5;
	wire bundleOut_0_a_valid = repeater_io_deq_valid;
	wire _T_8 = auto_out_a_ready & bundleOut_0_a_valid;
	wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 2'h0};
	wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1;
	wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1;
	wire [5:0] _GEN_9 = {4'd0, aFragOH1};
	wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_9;
	wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h03;
	wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4;
	wire [16:0] _GEN_10 = {11'd0, _bundleOut_0_a_bits_address_T_5};
	wire [3:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source, aToggle};
	wire _T_9 = ~repeater_io_full;
	TLMonitor_26 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	Repeater_6 repeater(
		.clock(repeater_clock),
		.reset(repeater_reset),
		.io_repeat(repeater_io_repeat),
		.io_full(repeater_io_full),
		.io_enq_ready(repeater_io_enq_ready),
		.io_enq_valid(repeater_io_enq_valid),
		.io_enq_bits_opcode(repeater_io_enq_bits_opcode),
		.io_enq_bits_param(repeater_io_enq_bits_param),
		.io_enq_bits_size(repeater_io_enq_bits_size),
		.io_enq_bits_source(repeater_io_enq_bits_source),
		.io_enq_bits_address(repeater_io_enq_bits_address),
		.io_enq_bits_mask(repeater_io_enq_bits_mask),
		.io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
		.io_deq_ready(repeater_io_deq_ready),
		.io_deq_valid(repeater_io_deq_valid),
		.io_deq_bits_opcode(repeater_io_deq_bits_opcode),
		.io_deq_bits_param(repeater_io_deq_bits_param),
		.io_deq_bits_size(repeater_io_deq_bits_size),
		.io_deq_bits_source(repeater_io_deq_bits_source),
		.io_deq_bits_address(repeater_io_deq_bits_address),
		.io_deq_bits_mask(repeater_io_deq_bits_mask),
		.io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = repeater_io_enq_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign auto_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_out_a_valid = repeater_io_deq_valid;
	assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode;
	assign auto_out_a_bits_param = repeater_io_deq_bits_param;
	assign auto_out_a_bits_size = aFrag[1:0];
	assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi, new_gennum};
	assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_10;
	assign auto_out_a_bits_mask = (repeater_io_full ? 4'hf : auto_in_a_bits_mask);
	assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = repeater_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid;
	assign monitor_io_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign repeater_clock = clock;
	assign repeater_reset = reset;
	assign repeater_io_repeat = new_gennum != 4'h0;
	assign repeater_io_enq_valid = auto_in_a_valid;
	assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign repeater_io_enq_bits_param = auto_in_a_bits_param;
	assign repeater_io_enq_bits_size = auto_in_a_bits_size;
	assign repeater_io_enq_bits_source = auto_in_a_bits_source;
	assign repeater_io_enq_bits_address = auto_in_a_bits_address;
	assign repeater_io_enq_bits_mask = auto_in_a_bits_mask;
	assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign repeater_io_deq_ready = auto_out_a_ready;
	always @(posedge clock) begin
		if (reset)
			acknum <= 4'h0;
		else if (_T_7)
			if (dFirst)
				acknum <= dFragnum;
			else
				acknum <= _acknum_T_1;
		if (_T_7)
			if (dFirst)
				dOrig <= dFirst_size;
		if (reset)
			dToggle <= 1'h0;
		else if (_T_7)
			if (dFirst)
				dToggle <= auto_out_d_bits_source[4];
		if (reset)
			gennum <= 4'h0;
		else if (_T_8)
			gennum <= new_gennum;
		if (aFirst)
			aToggle_r <= dToggle;
	end
endmodule
module TLInterconnectCoupler_14 (
	clock,
	reset,
	auto_fragmenter_out_a_ready,
	auto_fragmenter_out_a_valid,
	auto_fragmenter_out_a_bits_opcode,
	auto_fragmenter_out_a_bits_param,
	auto_fragmenter_out_a_bits_size,
	auto_fragmenter_out_a_bits_source,
	auto_fragmenter_out_a_bits_address,
	auto_fragmenter_out_a_bits_mask,
	auto_fragmenter_out_a_bits_corrupt,
	auto_fragmenter_out_d_ready,
	auto_fragmenter_out_d_valid,
	auto_fragmenter_out_d_bits_size,
	auto_fragmenter_out_d_bits_source,
	auto_fragmenter_out_d_bits_data,
	auto_tl_in_a_ready,
	auto_tl_in_a_valid,
	auto_tl_in_a_bits_opcode,
	auto_tl_in_a_bits_param,
	auto_tl_in_a_bits_size,
	auto_tl_in_a_bits_source,
	auto_tl_in_a_bits_address,
	auto_tl_in_a_bits_mask,
	auto_tl_in_a_bits_corrupt,
	auto_tl_in_d_ready,
	auto_tl_in_d_valid,
	auto_tl_in_d_bits_size,
	auto_tl_in_d_bits_source,
	auto_tl_in_d_bits_data
);
	input clock;
	input reset;
	input auto_fragmenter_out_a_ready;
	output wire auto_fragmenter_out_a_valid;
	output wire [2:0] auto_fragmenter_out_a_bits_opcode;
	output wire [2:0] auto_fragmenter_out_a_bits_param;
	output wire [1:0] auto_fragmenter_out_a_bits_size;
	output wire [7:0] auto_fragmenter_out_a_bits_source;
	output wire [16:0] auto_fragmenter_out_a_bits_address;
	output wire [3:0] auto_fragmenter_out_a_bits_mask;
	output wire auto_fragmenter_out_a_bits_corrupt;
	output wire auto_fragmenter_out_d_ready;
	input auto_fragmenter_out_d_valid;
	input [1:0] auto_fragmenter_out_d_bits_size;
	input [7:0] auto_fragmenter_out_d_bits_source;
	input [31:0] auto_fragmenter_out_d_bits_data;
	output wire auto_tl_in_a_ready;
	input auto_tl_in_a_valid;
	input [2:0] auto_tl_in_a_bits_opcode;
	input [2:0] auto_tl_in_a_bits_param;
	input [2:0] auto_tl_in_a_bits_size;
	input [2:0] auto_tl_in_a_bits_source;
	input [16:0] auto_tl_in_a_bits_address;
	input [3:0] auto_tl_in_a_bits_mask;
	input auto_tl_in_a_bits_corrupt;
	input auto_tl_in_d_ready;
	output wire auto_tl_in_d_valid;
	output wire [2:0] auto_tl_in_d_bits_size;
	output wire [2:0] auto_tl_in_d_bits_source;
	output wire [31:0] auto_tl_in_d_bits_data;
	wire fragmenter_clock;
	wire fragmenter_reset;
	wire fragmenter_auto_in_a_ready;
	wire fragmenter_auto_in_a_valid;
	wire [2:0] fragmenter_auto_in_a_bits_opcode;
	wire [2:0] fragmenter_auto_in_a_bits_param;
	wire [2:0] fragmenter_auto_in_a_bits_size;
	wire [2:0] fragmenter_auto_in_a_bits_source;
	wire [16:0] fragmenter_auto_in_a_bits_address;
	wire [3:0] fragmenter_auto_in_a_bits_mask;
	wire fragmenter_auto_in_a_bits_corrupt;
	wire fragmenter_auto_in_d_ready;
	wire fragmenter_auto_in_d_valid;
	wire [2:0] fragmenter_auto_in_d_bits_size;
	wire [2:0] fragmenter_auto_in_d_bits_source;
	wire [31:0] fragmenter_auto_in_d_bits_data;
	wire fragmenter_auto_out_a_ready;
	wire fragmenter_auto_out_a_valid;
	wire [2:0] fragmenter_auto_out_a_bits_opcode;
	wire [2:0] fragmenter_auto_out_a_bits_param;
	wire [1:0] fragmenter_auto_out_a_bits_size;
	wire [7:0] fragmenter_auto_out_a_bits_source;
	wire [16:0] fragmenter_auto_out_a_bits_address;
	wire [3:0] fragmenter_auto_out_a_bits_mask;
	wire fragmenter_auto_out_a_bits_corrupt;
	wire fragmenter_auto_out_d_ready;
	wire fragmenter_auto_out_d_valid;
	wire [1:0] fragmenter_auto_out_d_bits_size;
	wire [7:0] fragmenter_auto_out_d_bits_source;
	wire [31:0] fragmenter_auto_out_d_bits_data;
	TLFragmenter_5 fragmenter(
		.clock(fragmenter_clock),
		.reset(fragmenter_reset),
		.auto_in_a_ready(fragmenter_auto_in_a_ready),
		.auto_in_a_valid(fragmenter_auto_in_a_valid),
		.auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
		.auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
		.auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
		.auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
		.auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
		.auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
		.auto_in_d_ready(fragmenter_auto_in_d_ready),
		.auto_in_d_valid(fragmenter_auto_in_d_valid),
		.auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
		.auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
		.auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
		.auto_out_a_ready(fragmenter_auto_out_a_ready),
		.auto_out_a_valid(fragmenter_auto_out_a_valid),
		.auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
		.auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
		.auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
		.auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
		.auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
		.auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
		.auto_out_d_ready(fragmenter_auto_out_d_ready),
		.auto_out_d_valid(fragmenter_auto_out_d_valid),
		.auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
		.auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
		.auto_out_d_bits_data(fragmenter_auto_out_d_bits_data)
	);
	assign auto_fragmenter_out_a_valid = fragmenter_auto_out_a_valid;
	assign auto_fragmenter_out_a_bits_opcode = fragmenter_auto_out_a_bits_opcode;
	assign auto_fragmenter_out_a_bits_param = fragmenter_auto_out_a_bits_param;
	assign auto_fragmenter_out_a_bits_size = fragmenter_auto_out_a_bits_size;
	assign auto_fragmenter_out_a_bits_source = fragmenter_auto_out_a_bits_source;
	assign auto_fragmenter_out_a_bits_address = fragmenter_auto_out_a_bits_address;
	assign auto_fragmenter_out_a_bits_mask = fragmenter_auto_out_a_bits_mask;
	assign auto_fragmenter_out_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt;
	assign auto_fragmenter_out_d_ready = fragmenter_auto_out_d_ready;
	assign auto_tl_in_a_ready = fragmenter_auto_in_a_ready;
	assign auto_tl_in_d_valid = fragmenter_auto_in_d_valid;
	assign auto_tl_in_d_bits_size = fragmenter_auto_in_d_bits_size;
	assign auto_tl_in_d_bits_source = fragmenter_auto_in_d_bits_source;
	assign auto_tl_in_d_bits_data = fragmenter_auto_in_d_bits_data;
	assign fragmenter_clock = clock;
	assign fragmenter_reset = reset;
	assign fragmenter_auto_in_a_valid = auto_tl_in_a_valid;
	assign fragmenter_auto_in_a_bits_opcode = auto_tl_in_a_bits_opcode;
	assign fragmenter_auto_in_a_bits_param = auto_tl_in_a_bits_param;
	assign fragmenter_auto_in_a_bits_size = auto_tl_in_a_bits_size;
	assign fragmenter_auto_in_a_bits_source = auto_tl_in_a_bits_source;
	assign fragmenter_auto_in_a_bits_address = auto_tl_in_a_bits_address;
	assign fragmenter_auto_in_a_bits_mask = auto_tl_in_a_bits_mask;
	assign fragmenter_auto_in_a_bits_corrupt = auto_tl_in_a_bits_corrupt;
	assign fragmenter_auto_in_d_ready = auto_tl_in_d_ready;
	assign fragmenter_auto_out_a_ready = auto_fragmenter_out_a_ready;
	assign fragmenter_auto_out_d_valid = auto_fragmenter_out_d_valid;
	assign fragmenter_auto_out_d_bits_size = auto_fragmenter_out_d_bits_size;
	assign fragmenter_auto_out_d_bits_source = auto_fragmenter_out_d_bits_source;
	assign fragmenter_auto_out_d_bits_data = auto_fragmenter_out_d_bits_data;
endmodule
module TLInterconnectCoupler_15 (
	auto_tl_in_a_ready,
	auto_tl_in_a_valid,
	auto_tl_in_a_bits_address,
	auto_tl_in_a_bits_data,
	auto_tl_in_d_valid,
	auto_tl_out_a_ready,
	auto_tl_out_a_valid,
	auto_tl_out_a_bits_address,
	auto_tl_out_a_bits_data,
	auto_tl_out_d_valid
);
	output wire auto_tl_in_a_ready;
	input auto_tl_in_a_valid;
	input [31:0] auto_tl_in_a_bits_address;
	input [31:0] auto_tl_in_a_bits_data;
	output wire auto_tl_in_d_valid;
	input auto_tl_out_a_ready;
	output wire auto_tl_out_a_valid;
	output wire [31:0] auto_tl_out_a_bits_address;
	output wire [31:0] auto_tl_out_a_bits_data;
	input auto_tl_out_d_valid;
	assign auto_tl_in_a_ready = auto_tl_out_a_ready;
	assign auto_tl_in_d_valid = auto_tl_out_d_valid;
	assign auto_tl_out_a_valid = auto_tl_in_a_valid;
	assign auto_tl_out_a_bits_address = auto_tl_in_a_bits_address;
	assign auto_tl_out_a_bits_data = auto_tl_in_a_bits_data;
endmodule
module TLMonitor_27 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [1:0] io_in_a_bits_size;
	input [7:0] io_in_a_bits_source;
	input [20:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [1:0] io_in_d_bits_size;
	input [7:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_4 = io_in_a_bits_source <= 8'h9f;
	wire [4:0] _is_aligned_mask_T_1 = 5'h03 << io_in_a_bits_size;
	wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0];
	wire [20:0] _GEN_71 = {19'd0, is_aligned_mask};
	wire [20:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 21'h000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 2'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_10 = ~_source_ok_T_4;
	wire _T_20 = io_in_a_bits_opcode == 3'h6;
	wire [20:0] _T_33 = io_in_a_bits_address ^ 21'h100000;
	wire [21:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [21:0] _T_36 = $signed(_T_34) & -22'sh001000;
	wire _T_37 = $signed(_T_36) == 22'sh000000;
	wire _T_69 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_73 = ~io_in_a_bits_mask;
	wire _T_74 = _T_73 == 4'h0;
	wire _T_78 = ~io_in_a_bits_corrupt;
	wire _T_82 = io_in_a_bits_opcode == 3'h7;
	wire _T_135 = io_in_a_bits_param != 3'h0;
	wire _T_148 = io_in_a_bits_opcode == 3'h4;
	wire _T_164 = io_in_a_bits_size <= 2'h2;
	wire _T_172 = _T_164 & _T_37;
	wire _T_183 = io_in_a_bits_param == 3'h0;
	wire _T_187 = io_in_a_bits_mask == mask;
	wire _T_195 = io_in_a_bits_opcode == 3'h0;
	wire _T_218 = _source_ok_T_4 & _T_172;
	wire _T_236 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_273 = ~mask;
	wire [3:0] _T_274 = io_in_a_bits_mask & _T_273;
	wire _T_275 = _T_274 == 4'h0;
	wire _T_279 = io_in_a_bits_opcode == 3'h2;
	wire _T_309 = io_in_a_bits_param <= 3'h4;
	wire _T_317 = io_in_a_bits_opcode == 3'h3;
	wire _T_347 = io_in_a_bits_param <= 3'h3;
	wire _T_355 = io_in_a_bits_opcode == 3'h5;
	wire _T_385 = io_in_a_bits_param <= 3'h1;
	wire _T_397 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_10 = io_in_d_bits_source <= 8'h9f;
	wire _T_401 = io_in_d_bits_opcode == 3'h6;
	wire _T_405 = io_in_d_bits_size >= 2'h2;
	wire _T_409 = io_in_d_bits_param == 2'h0;
	wire _T_413 = ~io_in_d_bits_corrupt;
	wire _T_417 = ~io_in_d_bits_denied;
	wire _T_421 = io_in_d_bits_opcode == 3'h4;
	wire _T_432 = io_in_d_bits_param <= 2'h2;
	wire _T_436 = io_in_d_bits_param != 2'h2;
	wire _T_449 = io_in_d_bits_opcode == 3'h5;
	wire _T_469 = _T_417 | io_in_d_bits_corrupt;
	wire _T_478 = io_in_d_bits_opcode == 3'h0;
	wire _T_495 = io_in_d_bits_opcode == 3'h1;
	wire _T_513 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [1:0] size;
	reg [7:0] source;
	reg [20:0] address;
	wire _T_543 = io_in_a_valid & ~a_first;
	wire _T_544 = io_in_a_bits_opcode == opcode;
	wire _T_548 = io_in_a_bits_param == param;
	wire _T_552 = io_in_a_bits_size == size;
	wire _T_556 = io_in_a_bits_source == source;
	wire _T_560 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [1:0] size_1;
	reg [7:0] source_1;
	reg sink;
	reg denied;
	wire _T_567 = io_in_d_valid & ~d_first;
	wire _T_568 = io_in_d_bits_opcode == opcode_1;
	wire _T_572 = io_in_d_bits_param == param_1;
	wire _T_576 = io_in_d_bits_size == size_1;
	wire _T_580 = io_in_d_bits_source == source_1;
	wire _T_584 = io_in_d_bits_sink == sink;
	wire _T_588 = io_in_d_bits_denied == denied;
	reg [159:0] inflight;
	reg [639:0] inflight_opcodes;
	reg [639:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [10:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [639:0] _GEN_73 = {624'd0, _a_opcode_lookup_T_5};
	wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [639:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[639:1]};
	wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [639:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[639:1]};
	wire _T_594 = io_in_a_valid & a_first_1;
	wire [255:0] _a_set_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_a_bits_source;
	wire [255:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire _T_597 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1;
	wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [10:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [2050:0] _GEN_1 = {2047'd0, a_opcodes_set_interm};
	wire [2050:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? _a_sizes_set_interm_T_1 : 3'h0);
	wire [2049:0] _GEN_2 = {2047'd0, a_sizes_set_interm};
	wire [2049:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [159:0] _T_599 = inflight >> io_in_a_bits_source;
	wire _T_601 = ~_T_599[0];
	wire [255:0] _GEN_16 = (a_first_done & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2050:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 2051'h0);
	wire [2049:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 2050'h0);
	wire _T_605 = io_in_d_valid & d_first_1;
	wire _T_607 = ~_T_401;
	wire _T_608 = (io_in_d_valid & d_first_1) & ~_T_401;
	wire [255:0] _d_clr_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_d_bits_source;
	wire [255:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_401 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_3 = {2047'd0, _a_opcode_lookup_T_5};
	wire [2062:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [255:0] _GEN_22 = ((d_first_done & d_first_1) & _T_607 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_23 = ((d_first_done & d_first_1) & _T_607 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_594 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [159:0] _T_618 = inflight >> io_in_d_bits_source;
	wire _T_620 = _T_618[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_625 = io_in_d_bits_opcode == _GEN_40;
	wire _T_626 = (io_in_d_bits_opcode == _GEN_32) | _T_625;
	wire _T_630 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_637 = io_in_d_bits_opcode == _GEN_56;
	wire _T_638 = (io_in_d_bits_opcode == _GEN_48) | _T_637;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {2'd0, io_in_d_bits_size};
	wire _T_642 = _GEN_82 == a_size_lookup;
	wire _T_652 = (((_T_605 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_607;
	wire _T_654 = ~io_in_d_ready | io_in_a_ready;
	wire [159:0] a_set_wo_ready = _GEN_15[159:0];
	wire [159:0] d_clr_wo_ready = _GEN_21[159:0];
	wire _T_661 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [159:0] a_set = _GEN_16[159:0];
	wire [159:0] _inflight_T = inflight | a_set;
	wire [159:0] d_clr = _GEN_22[159:0];
	wire [159:0] _inflight_T_1 = ~d_clr;
	wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [639:0] a_opcodes_set = _GEN_19[639:0];
	wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [639:0] d_opcodes_clr = _GEN_23[639:0];
	wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [639:0] a_sizes_set = _GEN_20[639:0];
	wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_670 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [159:0] inflight_1;
	reg [639:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [639:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[639:1]};
	wire _T_696 = (io_in_d_valid & d_first_2) & _T_401;
	wire [255:0] _GEN_67 = ((d_first_done & d_first_2) & _T_401 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_68 = ((d_first_done & d_first_2) & _T_401 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire [159:0] _T_704 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_714 = _GEN_82 == c_size_lookup;
	wire [159:0] d_clr_1 = _GEN_67[159:0];
	wire [159:0] _inflight_T_4 = ~d_clr_1;
	wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0];
	wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_739 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			param <= io_in_a_bits_param;
		if (a_first_done & a_first)
			size <= io_in_a_bits_size;
		if (a_first_done & a_first)
			source <= io_in_a_bits_source;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			param_1 <= io_in_d_bits_param;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (d_first_done & d_first)
			sink <= io_in_d_bits_sink;
		if (d_first_done & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 160'h0000000000000000000000000000000000000000;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 640'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 640'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 160'h0000000000000000000000000000000000000000;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 640'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (d_first_done)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Queue_13 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_data,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [1:0] io_enq_bits_size;
	input [7:0] io_enq_bits_source;
	input [20:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input [31:0] io_enq_bits_data;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [1:0] io_deq_bits_size;
	output wire [7:0] io_deq_bits_source;
	output wire [20:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire [31:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg [2:0] ram_opcode [0:1];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [2:0] ram_param [0:1];
	wire ram_param_io_deq_bits_MPORT_en;
	wire ram_param_io_deq_bits_MPORT_addr;
	wire [2:0] ram_param_io_deq_bits_MPORT_data;
	wire [2:0] ram_param_MPORT_data;
	wire ram_param_MPORT_addr;
	wire ram_param_MPORT_mask;
	wire ram_param_MPORT_en;
	reg [1:0] ram_size [0:1];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [1:0] ram_size_io_deq_bits_MPORT_data;
	wire [1:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg [7:0] ram_source [0:1];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire [7:0] ram_source_io_deq_bits_MPORT_data;
	wire [7:0] ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg [20:0] ram_address [0:1];
	wire ram_address_io_deq_bits_MPORT_en;
	wire ram_address_io_deq_bits_MPORT_addr;
	wire [20:0] ram_address_io_deq_bits_MPORT_data;
	wire [20:0] ram_address_MPORT_data;
	wire ram_address_MPORT_addr;
	wire ram_address_MPORT_mask;
	wire ram_address_MPORT_en;
	reg [3:0] ram_mask [0:1];
	wire ram_mask_io_deq_bits_MPORT_en;
	wire ram_mask_io_deq_bits_MPORT_addr;
	wire [3:0] ram_mask_io_deq_bits_MPORT_data;
	wire [3:0] ram_mask_MPORT_data;
	wire ram_mask_MPORT_addr;
	wire ram_mask_MPORT_mask;
	wire ram_mask_MPORT_en;
	reg [31:0] ram_data [0:1];
	wire ram_data_io_deq_bits_MPORT_en;
	wire ram_data_io_deq_bits_MPORT_addr;
	wire [31:0] ram_data_io_deq_bits_MPORT_data;
	wire [31:0] ram_data_MPORT_data;
	wire ram_data_MPORT_addr;
	wire ram_data_MPORT_mask;
	wire ram_data_MPORT_en;
	reg ram_corrupt [0:1];
	wire ram_corrupt_io_deq_bits_MPORT_en;
	wire ram_corrupt_io_deq_bits_MPORT_addr;
	wire ram_corrupt_io_deq_bits_MPORT_data;
	wire ram_corrupt_MPORT_data;
	wire ram_corrupt_MPORT_addr;
	wire ram_corrupt_MPORT_mask;
	wire ram_corrupt_MPORT_en;
	reg value;
	reg value_1;
	reg maybe_full;
	wire ptr_match = value == value_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = value;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_param_io_deq_bits_MPORT_en = 1'h1;
	assign ram_param_io_deq_bits_MPORT_addr = value_1;
	assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr];
	assign ram_param_MPORT_data = io_enq_bits_param;
	assign ram_param_MPORT_addr = value;
	assign ram_param_MPORT_mask = 1'h1;
	assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = value_1;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = value;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = value_1;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = value;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_address_io_deq_bits_MPORT_en = 1'h1;
	assign ram_address_io_deq_bits_MPORT_addr = value_1;
	assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr];
	assign ram_address_MPORT_data = io_enq_bits_address;
	assign ram_address_MPORT_addr = value;
	assign ram_address_MPORT_mask = 1'h1;
	assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
	assign ram_mask_io_deq_bits_MPORT_addr = value_1;
	assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr];
	assign ram_mask_MPORT_data = io_enq_bits_mask;
	assign ram_mask_MPORT_addr = value;
	assign ram_mask_MPORT_mask = 1'h1;
	assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_data_io_deq_bits_MPORT_en = 1'h1;
	assign ram_data_io_deq_bits_MPORT_addr = value_1;
	assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr];
	assign ram_data_MPORT_data = io_enq_bits_data;
	assign ram_data_MPORT_addr = value;
	assign ram_data_MPORT_mask = 1'h1;
	assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
	assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
	assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr];
	assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
	assign ram_corrupt_MPORT_addr = value;
	assign ram_corrupt_MPORT_mask = 1'h1;
	assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data;
	assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data;
	assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data;
	assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_param_MPORT_en & ram_param_MPORT_mask)
			ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (ram_address_MPORT_en & ram_address_MPORT_mask)
			ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data;
		if (ram_mask_MPORT_en & ram_mask_MPORT_mask)
			ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data;
		if (ram_data_MPORT_en & ram_data_MPORT_mask)
			ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data;
		if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask)
			ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data;
		if (reset)
			value <= 1'h0;
		else if (do_enq)
			value <= value + 1'h1;
		if (reset)
			value_1 <= 1'h0;
		else if (do_deq)
			value_1 <= value_1 + 1'h1;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module Queue_14 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_data,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_sink,
	io_deq_bits_denied,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [1:0] io_enq_bits_size;
	input [7:0] io_enq_bits_source;
	input [31:0] io_enq_bits_data;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [1:0] io_deq_bits_param;
	output wire [1:0] io_deq_bits_size;
	output wire [7:0] io_deq_bits_source;
	output wire io_deq_bits_sink;
	output wire io_deq_bits_denied;
	output wire [31:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg [2:0] ram_opcode [0:1];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [1:0] ram_param [0:1];
	wire ram_param_io_deq_bits_MPORT_en;
	wire ram_param_io_deq_bits_MPORT_addr;
	wire [1:0] ram_param_io_deq_bits_MPORT_data;
	wire [1:0] ram_param_MPORT_data;
	wire ram_param_MPORT_addr;
	wire ram_param_MPORT_mask;
	wire ram_param_MPORT_en;
	reg [1:0] ram_size [0:1];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [1:0] ram_size_io_deq_bits_MPORT_data;
	wire [1:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg [7:0] ram_source [0:1];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire [7:0] ram_source_io_deq_bits_MPORT_data;
	wire [7:0] ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg ram_sink [0:1];
	wire ram_sink_io_deq_bits_MPORT_en;
	wire ram_sink_io_deq_bits_MPORT_addr;
	wire ram_sink_io_deq_bits_MPORT_data;
	wire ram_sink_MPORT_data;
	wire ram_sink_MPORT_addr;
	wire ram_sink_MPORT_mask;
	wire ram_sink_MPORT_en;
	reg ram_denied [0:1];
	wire ram_denied_io_deq_bits_MPORT_en;
	wire ram_denied_io_deq_bits_MPORT_addr;
	wire ram_denied_io_deq_bits_MPORT_data;
	wire ram_denied_MPORT_data;
	wire ram_denied_MPORT_addr;
	wire ram_denied_MPORT_mask;
	wire ram_denied_MPORT_en;
	reg [31:0] ram_data [0:1];
	wire ram_data_io_deq_bits_MPORT_en;
	wire ram_data_io_deq_bits_MPORT_addr;
	wire [31:0] ram_data_io_deq_bits_MPORT_data;
	wire [31:0] ram_data_MPORT_data;
	wire ram_data_MPORT_addr;
	wire ram_data_MPORT_mask;
	wire ram_data_MPORT_en;
	reg ram_corrupt [0:1];
	wire ram_corrupt_io_deq_bits_MPORT_en;
	wire ram_corrupt_io_deq_bits_MPORT_addr;
	wire ram_corrupt_io_deq_bits_MPORT_data;
	wire ram_corrupt_MPORT_data;
	wire ram_corrupt_MPORT_addr;
	wire ram_corrupt_MPORT_mask;
	wire ram_corrupt_MPORT_en;
	reg value;
	reg value_1;
	reg maybe_full;
	wire ptr_match = value == value_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = value;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_param_io_deq_bits_MPORT_en = 1'h1;
	assign ram_param_io_deq_bits_MPORT_addr = value_1;
	assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr];
	assign ram_param_MPORT_data = 2'h0;
	assign ram_param_MPORT_addr = value;
	assign ram_param_MPORT_mask = 1'h1;
	assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = value_1;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = value;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = value_1;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = value;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_sink_io_deq_bits_MPORT_en = 1'h1;
	assign ram_sink_io_deq_bits_MPORT_addr = value_1;
	assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr];
	assign ram_sink_MPORT_data = 1'h0;
	assign ram_sink_MPORT_addr = value;
	assign ram_sink_MPORT_mask = 1'h1;
	assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_denied_io_deq_bits_MPORT_en = 1'h1;
	assign ram_denied_io_deq_bits_MPORT_addr = value_1;
	assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr];
	assign ram_denied_MPORT_data = 1'h0;
	assign ram_denied_MPORT_addr = value;
	assign ram_denied_MPORT_mask = 1'h1;
	assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_data_io_deq_bits_MPORT_en = 1'h1;
	assign ram_data_io_deq_bits_MPORT_addr = value_1;
	assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr];
	assign ram_data_MPORT_data = io_enq_bits_data;
	assign ram_data_MPORT_addr = value;
	assign ram_data_MPORT_mask = 1'h1;
	assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
	assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
	assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr];
	assign ram_corrupt_MPORT_data = 1'h0;
	assign ram_corrupt_MPORT_addr = value;
	assign ram_corrupt_MPORT_mask = 1'h1;
	assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data;
	assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data;
	assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data;
	assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_param_MPORT_en & ram_param_MPORT_mask)
			ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (ram_sink_MPORT_en & ram_sink_MPORT_mask)
			ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data;
		if (ram_denied_MPORT_en & ram_denied_MPORT_mask)
			ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data;
		if (ram_data_MPORT_en & ram_data_MPORT_mask)
			ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data;
		if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask)
			ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data;
		if (reset)
			value <= 1'h0;
		else if (do_enq)
			value <= value + 1'h1;
		if (reset)
			value_1 <= 1'h0;
		else if (do_deq)
			value_1 <= value_1 + 1'h1;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module TLBuffer_9 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [1:0] auto_in_a_bits_size;
	input [7:0] auto_in_a_bits_source;
	input [20:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [1:0] auto_in_d_bits_size;
	output wire [7:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire [7:0] auto_out_a_bits_source;
	output wire [20:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_size;
	input [7:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [1:0] monitor_io_in_a_bits_size;
	wire [7:0] monitor_io_in_a_bits_source;
	wire [20:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [1:0] monitor_io_in_d_bits_size;
	wire [7:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire bundleOut_0_a_q_clock;
	wire bundleOut_0_a_q_reset;
	wire bundleOut_0_a_q_io_enq_ready;
	wire bundleOut_0_a_q_io_enq_valid;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_param;
	wire [1:0] bundleOut_0_a_q_io_enq_bits_size;
	wire [7:0] bundleOut_0_a_q_io_enq_bits_source;
	wire [20:0] bundleOut_0_a_q_io_enq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_data;
	wire bundleOut_0_a_q_io_enq_bits_corrupt;
	wire bundleOut_0_a_q_io_deq_ready;
	wire bundleOut_0_a_q_io_deq_valid;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_param;
	wire [1:0] bundleOut_0_a_q_io_deq_bits_size;
	wire [7:0] bundleOut_0_a_q_io_deq_bits_source;
	wire [20:0] bundleOut_0_a_q_io_deq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_data;
	wire bundleOut_0_a_q_io_deq_bits_corrupt;
	wire bundleIn_0_d_q_clock;
	wire bundleIn_0_d_q_reset;
	wire bundleIn_0_d_q_io_enq_ready;
	wire bundleIn_0_d_q_io_enq_valid;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_enq_bits_size;
	wire [7:0] bundleIn_0_d_q_io_enq_bits_source;
	wire [31:0] bundleIn_0_d_q_io_enq_bits_data;
	wire bundleIn_0_d_q_io_deq_ready;
	wire bundleIn_0_d_q_io_deq_valid;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_param;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_size;
	wire [7:0] bundleIn_0_d_q_io_deq_bits_source;
	wire bundleIn_0_d_q_io_deq_bits_sink;
	wire bundleIn_0_d_q_io_deq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_deq_bits_data;
	wire bundleIn_0_d_q_io_deq_bits_corrupt;
	TLMonitor_27 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Queue_13 bundleOut_0_a_q(
		.clock(bundleOut_0_a_q_clock),
		.reset(bundleOut_0_a_q_reset),
		.io_enq_ready(bundleOut_0_a_q_io_enq_ready),
		.io_enq_valid(bundleOut_0_a_q_io_enq_valid),
		.io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
		.io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
		.io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
		.io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
		.io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
		.io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleOut_0_a_q_io_deq_ready),
		.io_deq_valid(bundleOut_0_a_q_io_deq_valid),
		.io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
		.io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
		.io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
		.io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
		.io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
		.io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
	);
	Queue_14 bundleIn_0_d_q(
		.clock(bundleIn_0_d_q_clock),
		.reset(bundleIn_0_d_q_reset),
		.io_enq_ready(bundleIn_0_d_q_io_enq_ready),
		.io_enq_valid(bundleIn_0_d_q_io_enq_valid),
		.io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
		.io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
		.io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
		.io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
		.io_deq_ready(bundleIn_0_d_q_io_deq_ready),
		.io_deq_valid(bundleIn_0_d_q_io_deq_valid),
		.io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
		.io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
		.io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
		.io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
		.io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
		.io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data;
	assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid;
	assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode;
	assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param;
	assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size;
	assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source;
	assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address;
	assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask;
	assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data;
	assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt;
	assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign bundleOut_0_a_q_clock = clock;
	assign bundleOut_0_a_q_reset = reset;
	assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid;
	assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param;
	assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size;
	assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source;
	assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address;
	assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask;
	assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data;
	assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready;
	assign bundleIn_0_d_q_clock = clock;
	assign bundleIn_0_d_q_reset = reset;
	assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid;
	assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size;
	assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source;
	assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data;
	assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready;
endmodule
module TLMonitor_28 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [20:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [20:0] _GEN_71 = {15'd0, is_aligned_mask};
	wire [20:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 21'h000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [20:0] _T_56 = io_in_a_bits_address ^ 21'h100000;
	wire [21:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [21:0] _T_59 = $signed(_T_57) & -22'sh001000;
	wire _T_60 = $signed(_T_59) == 22'sh000000;
	wire _T_92 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_96 = ~io_in_a_bits_mask;
	wire _T_97 = _T_96 == 4'h0;
	wire _T_101 = ~io_in_a_bits_corrupt;
	wire _T_105 = io_in_a_bits_opcode == 3'h7;
	wire _T_159 = io_in_a_bits_param != 3'h0;
	wire _T_172 = io_in_a_bits_opcode == 3'h4;
	wire _T_189 = io_in_a_bits_size <= 3'h6;
	wire _T_197 = _T_189 & _T_60;
	wire _T_208 = io_in_a_bits_param == 3'h0;
	wire _T_212 = io_in_a_bits_mask == mask;
	wire _T_220 = io_in_a_bits_opcode == 3'h0;
	wire _T_244 = source_ok & _T_197;
	wire _T_262 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_300 = ~mask;
	wire [3:0] _T_301 = io_in_a_bits_mask & _T_300;
	wire _T_302 = _T_301 == 4'h0;
	wire _T_306 = io_in_a_bits_opcode == 3'h2;
	wire _T_337 = io_in_a_bits_param <= 3'h4;
	wire _T_345 = io_in_a_bits_opcode == 3'h3;
	wire _T_376 = io_in_a_bits_param <= 3'h3;
	wire _T_384 = io_in_a_bits_opcode == 3'h5;
	wire _T_415 = io_in_a_bits_param <= 3'h1;
	wire _T_427 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_431 = io_in_d_bits_opcode == 3'h6;
	wire _T_435 = io_in_d_bits_size >= 3'h2;
	wire _T_439 = io_in_d_bits_param == 2'h0;
	wire _T_443 = ~io_in_d_bits_corrupt;
	wire _T_447 = ~io_in_d_bits_denied;
	wire _T_451 = io_in_d_bits_opcode == 3'h4;
	wire _T_462 = io_in_d_bits_param <= 2'h2;
	wire _T_466 = io_in_d_bits_param != 2'h2;
	wire _T_479 = io_in_d_bits_opcode == 3'h5;
	wire _T_499 = _T_447 | io_in_d_bits_corrupt;
	wire _T_508 = io_in_d_bits_opcode == 3'h0;
	wire _T_525 = io_in_d_bits_opcode == 3'h1;
	wire _T_543 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [20:0] address;
	wire _T_573 = io_in_a_valid & ~a_first;
	wire _T_574 = io_in_a_bits_opcode == opcode;
	wire _T_578 = io_in_a_bits_param == param;
	wire _T_582 = io_in_a_bits_size == size;
	wire _T_586 = io_in_a_bits_source == source;
	wire _T_590 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_597 = io_in_d_valid & ~d_first;
	wire _T_598 = io_in_d_bits_opcode == opcode_1;
	wire _T_602 = io_in_d_bits_param == param_1;
	wire _T_606 = io_in_d_bits_size == size_1;
	wire _T_610 = io_in_d_bits_source == source_1;
	wire _T_614 = io_in_d_bits_sink == sink;
	wire _T_618 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_624 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire [7:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire _T_627 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_629 = inflight >> io_in_a_bits_source;
	wire _T_631 = ~_T_629[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_635 = io_in_d_valid & d_first_1;
	wire _T_637 = ~_T_431;
	wire _T_638 = (io_in_d_valid & d_first_1) & ~_T_431;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [7:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_431 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_637 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_637 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_624 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_648 = inflight >> io_in_d_bits_source;
	wire _T_650 = _T_648[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_655 = io_in_d_bits_opcode == _GEN_40;
	wire _T_656 = (io_in_d_bits_opcode == _GEN_32) | _T_655;
	wire _T_660 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_667 = io_in_d_bits_opcode == _GEN_56;
	wire _T_668 = (io_in_d_bits_opcode == _GEN_48) | _T_667;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_672 = _GEN_82 == a_size_lookup;
	wire _T_682 = (((_T_635 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_637;
	wire _T_684 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set_wo_ready = _GEN_15[4:0];
	wire [4:0] d_clr_wo_ready = _GEN_21[4:0];
	wire _T_691 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_700 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_726 = (io_in_d_valid & d_first_2) & _T_431;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_431 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_431 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_734 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_744 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_769 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Repeater_7 (
	clock,
	reset,
	io_repeat,
	io_full,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	input io_repeat;
	output wire io_full;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [20:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [20:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire io_deq_bits_corrupt;
	reg full;
	reg [2:0] saved_opcode;
	reg [2:0] saved_param;
	reg [2:0] saved_size;
	reg [2:0] saved_source;
	reg [20:0] saved_address;
	reg [3:0] saved_mask;
	reg saved_corrupt;
	wire _T = io_enq_ready & io_enq_valid;
	wire _GEN_0 = (_T & io_repeat) | full;
	wire _T_2 = io_deq_ready & io_deq_valid;
	assign io_full = full;
	assign io_enq_ready = io_deq_ready & ~full;
	assign io_deq_valid = io_enq_valid | full;
	assign io_deq_bits_opcode = (full ? saved_opcode : io_enq_bits_opcode);
	assign io_deq_bits_param = (full ? saved_param : io_enq_bits_param);
	assign io_deq_bits_size = (full ? saved_size : io_enq_bits_size);
	assign io_deq_bits_source = (full ? saved_source : io_enq_bits_source);
	assign io_deq_bits_address = (full ? saved_address : io_enq_bits_address);
	assign io_deq_bits_mask = (full ? saved_mask : io_enq_bits_mask);
	assign io_deq_bits_corrupt = (full ? saved_corrupt : io_enq_bits_corrupt);
	always @(posedge clock) begin
		if (reset)
			full <= 1'h0;
		else if (_T_2 & ~io_repeat)
			full <= 1'h0;
		else
			full <= _GEN_0;
		if (_T & io_repeat)
			saved_opcode <= io_enq_bits_opcode;
		if (_T & io_repeat)
			saved_param <= io_enq_bits_param;
		if (_T & io_repeat)
			saved_size <= io_enq_bits_size;
		if (_T & io_repeat)
			saved_source <= io_enq_bits_source;
		if (_T & io_repeat)
			saved_address <= io_enq_bits_address;
		if (_T & io_repeat)
			saved_mask <= io_enq_bits_mask;
		if (_T & io_repeat)
			saved_corrupt <= io_enq_bits_corrupt;
	end
endmodule
module TLFragmenter_6 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [20:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire [7:0] auto_out_a_bits_source;
	output wire [20:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [1:0] auto_out_d_bits_size;
	input [7:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [20:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire repeater_clock;
	wire repeater_reset;
	wire repeater_io_repeat;
	wire repeater_io_full;
	wire repeater_io_enq_ready;
	wire repeater_io_enq_valid;
	wire [2:0] repeater_io_enq_bits_opcode;
	wire [2:0] repeater_io_enq_bits_param;
	wire [2:0] repeater_io_enq_bits_size;
	wire [2:0] repeater_io_enq_bits_source;
	wire [20:0] repeater_io_enq_bits_address;
	wire [3:0] repeater_io_enq_bits_mask;
	wire repeater_io_enq_bits_corrupt;
	wire repeater_io_deq_ready;
	wire repeater_io_deq_valid;
	wire [2:0] repeater_io_deq_bits_opcode;
	wire [2:0] repeater_io_deq_bits_param;
	wire [2:0] repeater_io_deq_bits_size;
	wire [2:0] repeater_io_deq_bits_source;
	wire [20:0] repeater_io_deq_bits_address;
	wire [3:0] repeater_io_deq_bits_mask;
	wire repeater_io_deq_bits_corrupt;
	reg [3:0] acknum;
	reg [2:0] dOrig;
	reg dToggle;
	wire [3:0] dFragnum = auto_out_d_bits_source[3:0];
	wire dFirst = acknum == 4'h0;
	wire dLast = dFragnum == 4'h0;
	wire [3:0] _dsizeOH_T = 4'h1 << auto_out_d_bits_size;
	wire [2:0] dsizeOH = _dsizeOH_T[2:0];
	wire [4:0] _dsizeOH1_T_1 = 5'h03 << auto_out_d_bits_size;
	wire [1:0] dsizeOH1 = ~_dsizeOH1_T_1[1:0];
	wire dHasData = auto_out_d_bits_opcode[0];
	wire _T_5 = ~reset;
	wire ack_decrement = dHasData | dsizeOH[2];
	wire [5:0] _dFirst_size_T = {dFragnum, 2'h0};
	wire [5:0] _GEN_7 = {4'd0, dsizeOH1};
	wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7;
	wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0};
	wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h01;
	wire [6:0] _dFirst_size_T_4 = {1'h0, _dFirst_size_T_1};
	wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4;
	wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5;
	wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4];
	wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0];
	wire _dFirst_size_T_7 = |dFirst_size_hi;
	wire [3:0] _GEN_8 = {1'd0, dFirst_size_hi};
	wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo;
	wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2];
	wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0];
	wire _dFirst_size_T_9 = |dFirst_size_hi_1;
	wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1;
	wire [2:0] dFirst_size = {_dFirst_size_T_7, _dFirst_size_T_9, _dFirst_size_T_10[1]};
	wire drop = ~dHasData & ~dLast;
	wire bundleOut_0_d_ready = auto_in_d_ready | drop;
	wire _T_7 = bundleOut_0_d_ready & auto_out_d_valid;
	wire [3:0] _GEN_9 = {3'd0, ack_decrement};
	wire [3:0] _acknum_T_1 = acknum - _GEN_9;
	wire [2:0] aFrag = (repeater_io_deq_bits_size > 3'h2 ? 3'h2 : repeater_io_deq_bits_size);
	wire [12:0] _aOrigOH1_T_1 = 13'h003f << repeater_io_deq_bits_size;
	wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0];
	wire [8:0] _aFragOH1_T_1 = 9'h003 << aFrag;
	wire [1:0] aFragOH1 = ~_aFragOH1_T_1[1:0];
	wire aHasData = ~repeater_io_deq_bits_opcode[2];
	reg [3:0] gennum;
	wire aFirst = gennum == 4'h0;
	wire [3:0] _old_gennum1_T_2 = gennum - 4'h1;
	wire [3:0] old_gennum1 = (aFirst ? aOrigOH1[5:2] : _old_gennum1_T_2);
	wire [3:0] _new_gennum_T = ~old_gennum1;
	wire [3:0] new_gennum = ~_new_gennum_T;
	reg aToggle_r;
	wire _GEN_5 = (aFirst ? dToggle : aToggle_r);
	wire aToggle = ~_GEN_5;
	wire bundleOut_0_a_valid = repeater_io_deq_valid;
	wire _T_8 = auto_out_a_ready & bundleOut_0_a_valid;
	wire _repeater_io_repeat_T = ~aHasData;
	wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 2'h0};
	wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1;
	wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1;
	wire [5:0] _GEN_10 = {4'd0, aFragOH1};
	wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10;
	wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h03;
	wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4;
	wire [20:0] _GEN_11 = {15'd0, _bundleOut_0_a_bits_address_T_5};
	wire [3:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source, aToggle};
	wire _T_9 = ~repeater_io_full;
	TLMonitor_28 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Repeater_7 repeater(
		.clock(repeater_clock),
		.reset(repeater_reset),
		.io_repeat(repeater_io_repeat),
		.io_full(repeater_io_full),
		.io_enq_ready(repeater_io_enq_ready),
		.io_enq_valid(repeater_io_enq_valid),
		.io_enq_bits_opcode(repeater_io_enq_bits_opcode),
		.io_enq_bits_param(repeater_io_enq_bits_param),
		.io_enq_bits_size(repeater_io_enq_bits_size),
		.io_enq_bits_source(repeater_io_enq_bits_source),
		.io_enq_bits_address(repeater_io_enq_bits_address),
		.io_enq_bits_mask(repeater_io_enq_bits_mask),
		.io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
		.io_deq_ready(repeater_io_deq_ready),
		.io_deq_valid(repeater_io_deq_valid),
		.io_deq_bits_opcode(repeater_io_deq_bits_opcode),
		.io_deq_bits_param(repeater_io_deq_bits_param),
		.io_deq_bits_size(repeater_io_deq_bits_size),
		.io_deq_bits_source(repeater_io_deq_bits_source),
		.io_deq_bits_address(repeater_io_deq_bits_address),
		.io_deq_bits_mask(repeater_io_deq_bits_mask),
		.io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = repeater_io_enq_ready;
	assign auto_in_d_valid = auto_out_d_valid & ~drop;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign auto_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = repeater_io_deq_valid;
	assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode;
	assign auto_out_a_bits_param = repeater_io_deq_bits_param;
	assign auto_out_a_bits_size = aFrag[1:0];
	assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi, new_gennum};
	assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11;
	assign auto_out_a_bits_mask = (repeater_io_full ? 4'hf : auto_in_a_bits_mask);
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready | drop;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = repeater_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid & ~drop;
	assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_io_in_d_bits_param = auto_out_d_bits_param;
	assign monitor_io_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink;
	assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied;
	assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign repeater_clock = clock;
	assign repeater_reset = reset;
	assign repeater_io_repeat = ~aHasData & (new_gennum != 4'h0);
	assign repeater_io_enq_valid = auto_in_a_valid;
	assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign repeater_io_enq_bits_param = auto_in_a_bits_param;
	assign repeater_io_enq_bits_size = auto_in_a_bits_size;
	assign repeater_io_enq_bits_source = auto_in_a_bits_source;
	assign repeater_io_enq_bits_address = auto_in_a_bits_address;
	assign repeater_io_enq_bits_mask = auto_in_a_bits_mask;
	assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign repeater_io_deq_ready = auto_out_a_ready;
	always @(posedge clock) begin
		if (reset)
			acknum <= 4'h0;
		else if (_T_7)
			if (dFirst)
				acknum <= dFragnum;
			else
				acknum <= _acknum_T_1;
		if (_T_7)
			if (dFirst)
				dOrig <= dFirst_size;
		if (reset)
			dToggle <= 1'h0;
		else if (_T_7)
			if (dFirst)
				dToggle <= auto_out_d_bits_source[4];
		if (reset)
			gennum <= 4'h0;
		else if (_T_8)
			gennum <= new_gennum;
		if (aFirst)
			aToggle_r <= dToggle;
	end
endmodule
module TLBuffer_10 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [20:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [20:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module TLInterconnectCoupler_16 (
	clock,
	reset,
	auto_buffer_in_a_ready,
	auto_buffer_in_a_valid,
	auto_buffer_in_a_bits_opcode,
	auto_buffer_in_a_bits_param,
	auto_buffer_in_a_bits_size,
	auto_buffer_in_a_bits_source,
	auto_buffer_in_a_bits_address,
	auto_buffer_in_a_bits_mask,
	auto_buffer_in_a_bits_data,
	auto_buffer_in_a_bits_corrupt,
	auto_buffer_in_d_ready,
	auto_buffer_in_d_valid,
	auto_buffer_in_d_bits_opcode,
	auto_buffer_in_d_bits_param,
	auto_buffer_in_d_bits_size,
	auto_buffer_in_d_bits_source,
	auto_buffer_in_d_bits_sink,
	auto_buffer_in_d_bits_denied,
	auto_buffer_in_d_bits_data,
	auto_buffer_in_d_bits_corrupt,
	auto_buffer_out_a_ready,
	auto_buffer_out_a_valid,
	auto_buffer_out_a_bits_opcode,
	auto_buffer_out_a_bits_param,
	auto_buffer_out_a_bits_size,
	auto_buffer_out_a_bits_source,
	auto_buffer_out_a_bits_address,
	auto_buffer_out_a_bits_mask,
	auto_buffer_out_a_bits_data,
	auto_buffer_out_a_bits_corrupt,
	auto_buffer_out_d_ready,
	auto_buffer_out_d_valid,
	auto_buffer_out_d_bits_opcode,
	auto_buffer_out_d_bits_size,
	auto_buffer_out_d_bits_source,
	auto_buffer_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_buffer_in_a_ready;
	input auto_buffer_in_a_valid;
	input [2:0] auto_buffer_in_a_bits_opcode;
	input [2:0] auto_buffer_in_a_bits_param;
	input [2:0] auto_buffer_in_a_bits_size;
	input [2:0] auto_buffer_in_a_bits_source;
	input [20:0] auto_buffer_in_a_bits_address;
	input [3:0] auto_buffer_in_a_bits_mask;
	input [31:0] auto_buffer_in_a_bits_data;
	input auto_buffer_in_a_bits_corrupt;
	input auto_buffer_in_d_ready;
	output wire auto_buffer_in_d_valid;
	output wire [2:0] auto_buffer_in_d_bits_opcode;
	output wire [1:0] auto_buffer_in_d_bits_param;
	output wire [2:0] auto_buffer_in_d_bits_size;
	output wire [2:0] auto_buffer_in_d_bits_source;
	output wire auto_buffer_in_d_bits_sink;
	output wire auto_buffer_in_d_bits_denied;
	output wire [31:0] auto_buffer_in_d_bits_data;
	output wire auto_buffer_in_d_bits_corrupt;
	input auto_buffer_out_a_ready;
	output wire auto_buffer_out_a_valid;
	output wire [2:0] auto_buffer_out_a_bits_opcode;
	output wire [2:0] auto_buffer_out_a_bits_param;
	output wire [1:0] auto_buffer_out_a_bits_size;
	output wire [7:0] auto_buffer_out_a_bits_source;
	output wire [20:0] auto_buffer_out_a_bits_address;
	output wire [3:0] auto_buffer_out_a_bits_mask;
	output wire [31:0] auto_buffer_out_a_bits_data;
	output wire auto_buffer_out_a_bits_corrupt;
	output wire auto_buffer_out_d_ready;
	input auto_buffer_out_d_valid;
	input [2:0] auto_buffer_out_d_bits_opcode;
	input [1:0] auto_buffer_out_d_bits_size;
	input [7:0] auto_buffer_out_d_bits_source;
	input [31:0] auto_buffer_out_d_bits_data;
	wire buffer_clock;
	wire buffer_reset;
	wire buffer_auto_in_a_ready;
	wire buffer_auto_in_a_valid;
	wire [2:0] buffer_auto_in_a_bits_opcode;
	wire [2:0] buffer_auto_in_a_bits_param;
	wire [1:0] buffer_auto_in_a_bits_size;
	wire [7:0] buffer_auto_in_a_bits_source;
	wire [20:0] buffer_auto_in_a_bits_address;
	wire [3:0] buffer_auto_in_a_bits_mask;
	wire [31:0] buffer_auto_in_a_bits_data;
	wire buffer_auto_in_a_bits_corrupt;
	wire buffer_auto_in_d_ready;
	wire buffer_auto_in_d_valid;
	wire [2:0] buffer_auto_in_d_bits_opcode;
	wire [1:0] buffer_auto_in_d_bits_param;
	wire [1:0] buffer_auto_in_d_bits_size;
	wire [7:0] buffer_auto_in_d_bits_source;
	wire buffer_auto_in_d_bits_sink;
	wire buffer_auto_in_d_bits_denied;
	wire [31:0] buffer_auto_in_d_bits_data;
	wire buffer_auto_in_d_bits_corrupt;
	wire buffer_auto_out_a_ready;
	wire buffer_auto_out_a_valid;
	wire [2:0] buffer_auto_out_a_bits_opcode;
	wire [2:0] buffer_auto_out_a_bits_param;
	wire [1:0] buffer_auto_out_a_bits_size;
	wire [7:0] buffer_auto_out_a_bits_source;
	wire [20:0] buffer_auto_out_a_bits_address;
	wire [3:0] buffer_auto_out_a_bits_mask;
	wire [31:0] buffer_auto_out_a_bits_data;
	wire buffer_auto_out_a_bits_corrupt;
	wire buffer_auto_out_d_ready;
	wire buffer_auto_out_d_valid;
	wire [2:0] buffer_auto_out_d_bits_opcode;
	wire [1:0] buffer_auto_out_d_bits_size;
	wire [7:0] buffer_auto_out_d_bits_source;
	wire [31:0] buffer_auto_out_d_bits_data;
	wire fragmenter_clock;
	wire fragmenter_reset;
	wire fragmenter_auto_in_a_ready;
	wire fragmenter_auto_in_a_valid;
	wire [2:0] fragmenter_auto_in_a_bits_opcode;
	wire [2:0] fragmenter_auto_in_a_bits_param;
	wire [2:0] fragmenter_auto_in_a_bits_size;
	wire [2:0] fragmenter_auto_in_a_bits_source;
	wire [20:0] fragmenter_auto_in_a_bits_address;
	wire [3:0] fragmenter_auto_in_a_bits_mask;
	wire [31:0] fragmenter_auto_in_a_bits_data;
	wire fragmenter_auto_in_a_bits_corrupt;
	wire fragmenter_auto_in_d_ready;
	wire fragmenter_auto_in_d_valid;
	wire [2:0] fragmenter_auto_in_d_bits_opcode;
	wire [1:0] fragmenter_auto_in_d_bits_param;
	wire [2:0] fragmenter_auto_in_d_bits_size;
	wire [2:0] fragmenter_auto_in_d_bits_source;
	wire fragmenter_auto_in_d_bits_sink;
	wire fragmenter_auto_in_d_bits_denied;
	wire [31:0] fragmenter_auto_in_d_bits_data;
	wire fragmenter_auto_in_d_bits_corrupt;
	wire fragmenter_auto_out_a_ready;
	wire fragmenter_auto_out_a_valid;
	wire [2:0] fragmenter_auto_out_a_bits_opcode;
	wire [2:0] fragmenter_auto_out_a_bits_param;
	wire [1:0] fragmenter_auto_out_a_bits_size;
	wire [7:0] fragmenter_auto_out_a_bits_source;
	wire [20:0] fragmenter_auto_out_a_bits_address;
	wire [3:0] fragmenter_auto_out_a_bits_mask;
	wire [31:0] fragmenter_auto_out_a_bits_data;
	wire fragmenter_auto_out_a_bits_corrupt;
	wire fragmenter_auto_out_d_ready;
	wire fragmenter_auto_out_d_valid;
	wire [2:0] fragmenter_auto_out_d_bits_opcode;
	wire [1:0] fragmenter_auto_out_d_bits_param;
	wire [1:0] fragmenter_auto_out_d_bits_size;
	wire [7:0] fragmenter_auto_out_d_bits_source;
	wire fragmenter_auto_out_d_bits_sink;
	wire fragmenter_auto_out_d_bits_denied;
	wire [31:0] fragmenter_auto_out_d_bits_data;
	wire fragmenter_auto_out_d_bits_corrupt;
	wire buffer_1_auto_in_a_ready;
	wire buffer_1_auto_in_a_valid;
	wire [2:0] buffer_1_auto_in_a_bits_opcode;
	wire [2:0] buffer_1_auto_in_a_bits_param;
	wire [2:0] buffer_1_auto_in_a_bits_size;
	wire [2:0] buffer_1_auto_in_a_bits_source;
	wire [20:0] buffer_1_auto_in_a_bits_address;
	wire [3:0] buffer_1_auto_in_a_bits_mask;
	wire [31:0] buffer_1_auto_in_a_bits_data;
	wire buffer_1_auto_in_a_bits_corrupt;
	wire buffer_1_auto_in_d_ready;
	wire buffer_1_auto_in_d_valid;
	wire [2:0] buffer_1_auto_in_d_bits_opcode;
	wire [1:0] buffer_1_auto_in_d_bits_param;
	wire [2:0] buffer_1_auto_in_d_bits_size;
	wire [2:0] buffer_1_auto_in_d_bits_source;
	wire buffer_1_auto_in_d_bits_sink;
	wire buffer_1_auto_in_d_bits_denied;
	wire [31:0] buffer_1_auto_in_d_bits_data;
	wire buffer_1_auto_in_d_bits_corrupt;
	wire buffer_1_auto_out_a_ready;
	wire buffer_1_auto_out_a_valid;
	wire [2:0] buffer_1_auto_out_a_bits_opcode;
	wire [2:0] buffer_1_auto_out_a_bits_param;
	wire [2:0] buffer_1_auto_out_a_bits_size;
	wire [2:0] buffer_1_auto_out_a_bits_source;
	wire [20:0] buffer_1_auto_out_a_bits_address;
	wire [3:0] buffer_1_auto_out_a_bits_mask;
	wire [31:0] buffer_1_auto_out_a_bits_data;
	wire buffer_1_auto_out_a_bits_corrupt;
	wire buffer_1_auto_out_d_ready;
	wire buffer_1_auto_out_d_valid;
	wire [2:0] buffer_1_auto_out_d_bits_opcode;
	wire [1:0] buffer_1_auto_out_d_bits_param;
	wire [2:0] buffer_1_auto_out_d_bits_size;
	wire [2:0] buffer_1_auto_out_d_bits_source;
	wire buffer_1_auto_out_d_bits_sink;
	wire buffer_1_auto_out_d_bits_denied;
	wire [31:0] buffer_1_auto_out_d_bits_data;
	wire buffer_1_auto_out_d_bits_corrupt;
	TLBuffer_9 buffer(
		.clock(buffer_clock),
		.reset(buffer_reset),
		.auto_in_a_ready(buffer_auto_in_a_ready),
		.auto_in_a_valid(buffer_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_auto_in_d_ready),
		.auto_in_d_valid(buffer_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_auto_out_a_ready),
		.auto_out_a_valid(buffer_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_auto_out_d_ready),
		.auto_out_d_valid(buffer_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(buffer_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_auto_out_d_bits_source),
		.auto_out_d_bits_data(buffer_auto_out_d_bits_data)
	);
	TLFragmenter_6 fragmenter(
		.clock(fragmenter_clock),
		.reset(fragmenter_reset),
		.auto_in_a_ready(fragmenter_auto_in_a_ready),
		.auto_in_a_valid(fragmenter_auto_in_a_valid),
		.auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
		.auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
		.auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
		.auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
		.auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
		.auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
		.auto_in_d_ready(fragmenter_auto_in_d_ready),
		.auto_in_d_valid(fragmenter_auto_in_d_valid),
		.auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(fragmenter_auto_in_d_bits_param),
		.auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
		.auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
		.auto_in_d_bits_sink(fragmenter_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(fragmenter_auto_in_d_bits_denied),
		.auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(fragmenter_auto_in_d_bits_corrupt),
		.auto_out_a_ready(fragmenter_auto_out_a_ready),
		.auto_out_a_valid(fragmenter_auto_out_a_valid),
		.auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
		.auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
		.auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
		.auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
		.auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
		.auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
		.auto_out_d_ready(fragmenter_auto_out_d_ready),
		.auto_out_d_valid(fragmenter_auto_out_d_valid),
		.auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(fragmenter_auto_out_d_bits_param),
		.auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
		.auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
		.auto_out_d_bits_sink(fragmenter_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(fragmenter_auto_out_d_bits_denied),
		.auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(fragmenter_auto_out_d_bits_corrupt)
	);
	TLBuffer_10 buffer_1(
		.auto_in_a_ready(buffer_1_auto_in_a_ready),
		.auto_in_a_valid(buffer_1_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_1_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_1_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_1_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_1_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_1_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_1_auto_in_d_ready),
		.auto_in_d_valid(buffer_1_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_1_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_1_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_1_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_1_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_1_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_1_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_1_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_1_auto_out_a_ready),
		.auto_out_a_valid(buffer_1_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_1_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_1_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_1_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_1_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_1_auto_out_d_ready),
		.auto_out_d_valid(buffer_1_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(buffer_1_auto_out_d_bits_param),
		.auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
		.auto_out_d_bits_sink(buffer_1_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
		.auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt)
	);
	assign auto_buffer_in_a_ready = buffer_1_auto_in_a_ready;
	assign auto_buffer_in_d_valid = buffer_1_auto_in_d_valid;
	assign auto_buffer_in_d_bits_opcode = buffer_1_auto_in_d_bits_opcode;
	assign auto_buffer_in_d_bits_param = buffer_1_auto_in_d_bits_param;
	assign auto_buffer_in_d_bits_size = buffer_1_auto_in_d_bits_size;
	assign auto_buffer_in_d_bits_source = buffer_1_auto_in_d_bits_source;
	assign auto_buffer_in_d_bits_sink = buffer_1_auto_in_d_bits_sink;
	assign auto_buffer_in_d_bits_denied = buffer_1_auto_in_d_bits_denied;
	assign auto_buffer_in_d_bits_data = buffer_1_auto_in_d_bits_data;
	assign auto_buffer_in_d_bits_corrupt = buffer_1_auto_in_d_bits_corrupt;
	assign auto_buffer_out_a_valid = buffer_auto_out_a_valid;
	assign auto_buffer_out_a_bits_opcode = buffer_auto_out_a_bits_opcode;
	assign auto_buffer_out_a_bits_param = buffer_auto_out_a_bits_param;
	assign auto_buffer_out_a_bits_size = buffer_auto_out_a_bits_size;
	assign auto_buffer_out_a_bits_source = buffer_auto_out_a_bits_source;
	assign auto_buffer_out_a_bits_address = buffer_auto_out_a_bits_address;
	assign auto_buffer_out_a_bits_mask = buffer_auto_out_a_bits_mask;
	assign auto_buffer_out_a_bits_data = buffer_auto_out_a_bits_data;
	assign auto_buffer_out_a_bits_corrupt = buffer_auto_out_a_bits_corrupt;
	assign auto_buffer_out_d_ready = buffer_auto_out_d_ready;
	assign buffer_clock = clock;
	assign buffer_reset = reset;
	assign buffer_auto_in_a_valid = fragmenter_auto_out_a_valid;
	assign buffer_auto_in_a_bits_opcode = fragmenter_auto_out_a_bits_opcode;
	assign buffer_auto_in_a_bits_param = fragmenter_auto_out_a_bits_param;
	assign buffer_auto_in_a_bits_size = fragmenter_auto_out_a_bits_size;
	assign buffer_auto_in_a_bits_source = fragmenter_auto_out_a_bits_source;
	assign buffer_auto_in_a_bits_address = fragmenter_auto_out_a_bits_address;
	assign buffer_auto_in_a_bits_mask = fragmenter_auto_out_a_bits_mask;
	assign buffer_auto_in_a_bits_data = fragmenter_auto_out_a_bits_data;
	assign buffer_auto_in_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt;
	assign buffer_auto_in_d_ready = fragmenter_auto_out_d_ready;
	assign buffer_auto_out_a_ready = auto_buffer_out_a_ready;
	assign buffer_auto_out_d_valid = auto_buffer_out_d_valid;
	assign buffer_auto_out_d_bits_opcode = auto_buffer_out_d_bits_opcode;
	assign buffer_auto_out_d_bits_size = auto_buffer_out_d_bits_size;
	assign buffer_auto_out_d_bits_source = auto_buffer_out_d_bits_source;
	assign buffer_auto_out_d_bits_data = auto_buffer_out_d_bits_data;
	assign fragmenter_clock = clock;
	assign fragmenter_reset = reset;
	assign fragmenter_auto_in_a_valid = buffer_1_auto_out_a_valid;
	assign fragmenter_auto_in_a_bits_opcode = buffer_1_auto_out_a_bits_opcode;
	assign fragmenter_auto_in_a_bits_param = buffer_1_auto_out_a_bits_param;
	assign fragmenter_auto_in_a_bits_size = buffer_1_auto_out_a_bits_size;
	assign fragmenter_auto_in_a_bits_source = buffer_1_auto_out_a_bits_source;
	assign fragmenter_auto_in_a_bits_address = buffer_1_auto_out_a_bits_address;
	assign fragmenter_auto_in_a_bits_mask = buffer_1_auto_out_a_bits_mask;
	assign fragmenter_auto_in_a_bits_data = buffer_1_auto_out_a_bits_data;
	assign fragmenter_auto_in_a_bits_corrupt = buffer_1_auto_out_a_bits_corrupt;
	assign fragmenter_auto_in_d_ready = buffer_1_auto_out_d_ready;
	assign fragmenter_auto_out_a_ready = buffer_auto_in_a_ready;
	assign fragmenter_auto_out_d_valid = buffer_auto_in_d_valid;
	assign fragmenter_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode;
	assign fragmenter_auto_out_d_bits_param = buffer_auto_in_d_bits_param;
	assign fragmenter_auto_out_d_bits_size = buffer_auto_in_d_bits_size;
	assign fragmenter_auto_out_d_bits_source = buffer_auto_in_d_bits_source;
	assign fragmenter_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink;
	assign fragmenter_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied;
	assign fragmenter_auto_out_d_bits_data = buffer_auto_in_d_bits_data;
	assign fragmenter_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt;
	assign buffer_1_auto_in_a_valid = auto_buffer_in_a_valid;
	assign buffer_1_auto_in_a_bits_opcode = auto_buffer_in_a_bits_opcode;
	assign buffer_1_auto_in_a_bits_param = auto_buffer_in_a_bits_param;
	assign buffer_1_auto_in_a_bits_size = auto_buffer_in_a_bits_size;
	assign buffer_1_auto_in_a_bits_source = auto_buffer_in_a_bits_source;
	assign buffer_1_auto_in_a_bits_address = auto_buffer_in_a_bits_address;
	assign buffer_1_auto_in_a_bits_mask = auto_buffer_in_a_bits_mask;
	assign buffer_1_auto_in_a_bits_data = auto_buffer_in_a_bits_data;
	assign buffer_1_auto_in_a_bits_corrupt = auto_buffer_in_a_bits_corrupt;
	assign buffer_1_auto_in_d_ready = auto_buffer_in_d_ready;
	assign buffer_1_auto_out_a_ready = fragmenter_auto_in_a_ready;
	assign buffer_1_auto_out_d_valid = fragmenter_auto_in_d_valid;
	assign buffer_1_auto_out_d_bits_opcode = fragmenter_auto_in_d_bits_opcode;
	assign buffer_1_auto_out_d_bits_param = fragmenter_auto_in_d_bits_param;
	assign buffer_1_auto_out_d_bits_size = fragmenter_auto_in_d_bits_size;
	assign buffer_1_auto_out_d_bits_source = fragmenter_auto_in_d_bits_source;
	assign buffer_1_auto_out_d_bits_sink = fragmenter_auto_in_d_bits_sink;
	assign buffer_1_auto_out_d_bits_denied = fragmenter_auto_in_d_bits_denied;
	assign buffer_1_auto_out_d_bits_data = fragmenter_auto_in_d_bits_data;
	assign buffer_1_auto_out_d_bits_corrupt = fragmenter_auto_in_d_bits_corrupt;
endmodule
module TLMonitor_29 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [1:0] io_in_a_bits_size;
	input [7:0] io_in_a_bits_source;
	input [20:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [1:0] io_in_d_bits_size;
	input [7:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_4 = io_in_a_bits_source <= 8'h9f;
	wire [4:0] _is_aligned_mask_T_1 = 5'h03 << io_in_a_bits_size;
	wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0];
	wire [20:0] _GEN_71 = {19'd0, is_aligned_mask};
	wire [20:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 21'h000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 2'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_10 = ~_source_ok_T_4;
	wire _T_20 = io_in_a_bits_opcode == 3'h6;
	wire [20:0] _T_33 = io_in_a_bits_address ^ 21'h110000;
	wire [21:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [21:0] _T_36 = $signed(_T_34) & -22'sh001000;
	wire _T_37 = $signed(_T_36) == 22'sh000000;
	wire _T_69 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_73 = ~io_in_a_bits_mask;
	wire _T_74 = _T_73 == 4'h0;
	wire _T_78 = ~io_in_a_bits_corrupt;
	wire _T_82 = io_in_a_bits_opcode == 3'h7;
	wire _T_135 = io_in_a_bits_param != 3'h0;
	wire _T_148 = io_in_a_bits_opcode == 3'h4;
	wire _T_164 = io_in_a_bits_size <= 2'h2;
	wire _T_172 = _T_164 & _T_37;
	wire _T_183 = io_in_a_bits_param == 3'h0;
	wire _T_187 = io_in_a_bits_mask == mask;
	wire _T_195 = io_in_a_bits_opcode == 3'h0;
	wire _T_218 = _source_ok_T_4 & _T_172;
	wire _T_236 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_273 = ~mask;
	wire [3:0] _T_274 = io_in_a_bits_mask & _T_273;
	wire _T_275 = _T_274 == 4'h0;
	wire _T_279 = io_in_a_bits_opcode == 3'h2;
	wire _T_309 = io_in_a_bits_param <= 3'h4;
	wire _T_317 = io_in_a_bits_opcode == 3'h3;
	wire _T_347 = io_in_a_bits_param <= 3'h3;
	wire _T_355 = io_in_a_bits_opcode == 3'h5;
	wire _T_385 = io_in_a_bits_param <= 3'h1;
	wire _T_397 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_10 = io_in_d_bits_source <= 8'h9f;
	wire _T_401 = io_in_d_bits_opcode == 3'h6;
	wire _T_405 = io_in_d_bits_size >= 2'h2;
	wire _T_409 = io_in_d_bits_param == 2'h0;
	wire _T_413 = ~io_in_d_bits_corrupt;
	wire _T_417 = ~io_in_d_bits_denied;
	wire _T_421 = io_in_d_bits_opcode == 3'h4;
	wire _T_432 = io_in_d_bits_param <= 2'h2;
	wire _T_436 = io_in_d_bits_param != 2'h2;
	wire _T_449 = io_in_d_bits_opcode == 3'h5;
	wire _T_469 = _T_417 | io_in_d_bits_corrupt;
	wire _T_478 = io_in_d_bits_opcode == 3'h0;
	wire _T_495 = io_in_d_bits_opcode == 3'h1;
	wire _T_513 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [1:0] size;
	reg [7:0] source;
	reg [20:0] address;
	wire _T_543 = io_in_a_valid & ~a_first;
	wire _T_544 = io_in_a_bits_opcode == opcode;
	wire _T_548 = io_in_a_bits_param == param;
	wire _T_552 = io_in_a_bits_size == size;
	wire _T_556 = io_in_a_bits_source == source;
	wire _T_560 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [1:0] size_1;
	reg [7:0] source_1;
	reg sink;
	reg denied;
	wire _T_567 = io_in_d_valid & ~d_first;
	wire _T_568 = io_in_d_bits_opcode == opcode_1;
	wire _T_572 = io_in_d_bits_param == param_1;
	wire _T_576 = io_in_d_bits_size == size_1;
	wire _T_580 = io_in_d_bits_source == source_1;
	wire _T_584 = io_in_d_bits_sink == sink;
	wire _T_588 = io_in_d_bits_denied == denied;
	reg [159:0] inflight;
	reg [639:0] inflight_opcodes;
	reg [639:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [10:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [639:0] _GEN_73 = {624'd0, _a_opcode_lookup_T_5};
	wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [639:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[639:1]};
	wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [639:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[639:1]};
	wire _T_594 = io_in_a_valid & a_first_1;
	wire [255:0] _a_set_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_a_bits_source;
	wire [255:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire _T_597 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1;
	wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [10:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [2050:0] _GEN_1 = {2047'd0, a_opcodes_set_interm};
	wire [2050:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? _a_sizes_set_interm_T_1 : 3'h0);
	wire [2049:0] _GEN_2 = {2047'd0, a_sizes_set_interm};
	wire [2049:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [159:0] _T_599 = inflight >> io_in_a_bits_source;
	wire _T_601 = ~_T_599[0];
	wire [255:0] _GEN_16 = (a_first_done & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2050:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 2051'h0);
	wire [2049:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 2050'h0);
	wire _T_605 = io_in_d_valid & d_first_1;
	wire _T_607 = ~_T_401;
	wire _T_608 = (io_in_d_valid & d_first_1) & ~_T_401;
	wire [255:0] _d_clr_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_d_bits_source;
	wire [255:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_401 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_3 = {2047'd0, _a_opcode_lookup_T_5};
	wire [2062:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [255:0] _GEN_22 = ((d_first_done & d_first_1) & _T_607 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_23 = ((d_first_done & d_first_1) & _T_607 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_594 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [159:0] _T_618 = inflight >> io_in_d_bits_source;
	wire _T_620 = _T_618[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_625 = io_in_d_bits_opcode == _GEN_40;
	wire _T_626 = (io_in_d_bits_opcode == _GEN_32) | _T_625;
	wire _T_630 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_637 = io_in_d_bits_opcode == _GEN_56;
	wire _T_638 = (io_in_d_bits_opcode == _GEN_48) | _T_637;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {2'd0, io_in_d_bits_size};
	wire _T_642 = _GEN_82 == a_size_lookup;
	wire _T_652 = (((_T_605 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_607;
	wire _T_654 = ~io_in_d_ready | io_in_a_ready;
	wire [159:0] a_set_wo_ready = _GEN_15[159:0];
	wire [159:0] d_clr_wo_ready = _GEN_21[159:0];
	wire _T_661 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [159:0] a_set = _GEN_16[159:0];
	wire [159:0] _inflight_T = inflight | a_set;
	wire [159:0] d_clr = _GEN_22[159:0];
	wire [159:0] _inflight_T_1 = ~d_clr;
	wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [639:0] a_opcodes_set = _GEN_19[639:0];
	wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [639:0] d_opcodes_clr = _GEN_23[639:0];
	wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [639:0] a_sizes_set = _GEN_20[639:0];
	wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_670 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [159:0] inflight_1;
	reg [639:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [639:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[639:1]};
	wire _T_696 = (io_in_d_valid & d_first_2) & _T_401;
	wire [255:0] _GEN_67 = ((d_first_done & d_first_2) & _T_401 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_68 = ((d_first_done & d_first_2) & _T_401 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire [159:0] _T_704 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_714 = _GEN_82 == c_size_lookup;
	wire [159:0] d_clr_1 = _GEN_67[159:0];
	wire [159:0] _inflight_T_4 = ~d_clr_1;
	wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0];
	wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_739 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			param <= io_in_a_bits_param;
		if (a_first_done & a_first)
			size <= io_in_a_bits_size;
		if (a_first_done & a_first)
			source <= io_in_a_bits_source;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			param_1 <= io_in_d_bits_param;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (d_first_done & d_first)
			sink <= io_in_d_bits_sink;
		if (d_first_done & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 160'h0000000000000000000000000000000000000000;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 640'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 640'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 160'h0000000000000000000000000000000000000000;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 640'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (d_first_done)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLBuffer_11 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [1:0] auto_in_a_bits_size;
	input [7:0] auto_in_a_bits_source;
	input [20:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [1:0] auto_in_d_bits_size;
	output wire [7:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire [7:0] auto_out_a_bits_source;
	output wire [20:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_size;
	input [7:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [1:0] monitor_io_in_a_bits_size;
	wire [7:0] monitor_io_in_a_bits_source;
	wire [20:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [1:0] monitor_io_in_d_bits_size;
	wire [7:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire bundleOut_0_a_q_clock;
	wire bundleOut_0_a_q_reset;
	wire bundleOut_0_a_q_io_enq_ready;
	wire bundleOut_0_a_q_io_enq_valid;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_param;
	wire [1:0] bundleOut_0_a_q_io_enq_bits_size;
	wire [7:0] bundleOut_0_a_q_io_enq_bits_source;
	wire [20:0] bundleOut_0_a_q_io_enq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_data;
	wire bundleOut_0_a_q_io_enq_bits_corrupt;
	wire bundleOut_0_a_q_io_deq_ready;
	wire bundleOut_0_a_q_io_deq_valid;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_param;
	wire [1:0] bundleOut_0_a_q_io_deq_bits_size;
	wire [7:0] bundleOut_0_a_q_io_deq_bits_source;
	wire [20:0] bundleOut_0_a_q_io_deq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_data;
	wire bundleOut_0_a_q_io_deq_bits_corrupt;
	wire bundleIn_0_d_q_clock;
	wire bundleIn_0_d_q_reset;
	wire bundleIn_0_d_q_io_enq_ready;
	wire bundleIn_0_d_q_io_enq_valid;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_enq_bits_size;
	wire [7:0] bundleIn_0_d_q_io_enq_bits_source;
	wire [31:0] bundleIn_0_d_q_io_enq_bits_data;
	wire bundleIn_0_d_q_io_deq_ready;
	wire bundleIn_0_d_q_io_deq_valid;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_param;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_size;
	wire [7:0] bundleIn_0_d_q_io_deq_bits_source;
	wire bundleIn_0_d_q_io_deq_bits_sink;
	wire bundleIn_0_d_q_io_deq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_deq_bits_data;
	wire bundleIn_0_d_q_io_deq_bits_corrupt;
	TLMonitor_29 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Queue_13 bundleOut_0_a_q(
		.clock(bundleOut_0_a_q_clock),
		.reset(bundleOut_0_a_q_reset),
		.io_enq_ready(bundleOut_0_a_q_io_enq_ready),
		.io_enq_valid(bundleOut_0_a_q_io_enq_valid),
		.io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
		.io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
		.io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
		.io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
		.io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
		.io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleOut_0_a_q_io_deq_ready),
		.io_deq_valid(bundleOut_0_a_q_io_deq_valid),
		.io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
		.io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
		.io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
		.io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
		.io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
		.io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
	);
	Queue_14 bundleIn_0_d_q(
		.clock(bundleIn_0_d_q_clock),
		.reset(bundleIn_0_d_q_reset),
		.io_enq_ready(bundleIn_0_d_q_io_enq_ready),
		.io_enq_valid(bundleIn_0_d_q_io_enq_valid),
		.io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
		.io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
		.io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
		.io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
		.io_deq_ready(bundleIn_0_d_q_io_deq_ready),
		.io_deq_valid(bundleIn_0_d_q_io_deq_valid),
		.io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
		.io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
		.io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
		.io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
		.io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
		.io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data;
	assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid;
	assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode;
	assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param;
	assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size;
	assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source;
	assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address;
	assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask;
	assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data;
	assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt;
	assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign bundleOut_0_a_q_clock = clock;
	assign bundleOut_0_a_q_reset = reset;
	assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid;
	assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param;
	assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size;
	assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source;
	assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address;
	assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask;
	assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data;
	assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready;
	assign bundleIn_0_d_q_clock = clock;
	assign bundleIn_0_d_q_reset = reset;
	assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid;
	assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size;
	assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source;
	assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data;
	assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready;
endmodule
module TLMonitor_30 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [20:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [20:0] _GEN_71 = {15'd0, is_aligned_mask};
	wire [20:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 21'h000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [20:0] _T_56 = io_in_a_bits_address ^ 21'h110000;
	wire [21:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [21:0] _T_59 = $signed(_T_57) & -22'sh001000;
	wire _T_60 = $signed(_T_59) == 22'sh000000;
	wire _T_92 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_96 = ~io_in_a_bits_mask;
	wire _T_97 = _T_96 == 4'h0;
	wire _T_101 = ~io_in_a_bits_corrupt;
	wire _T_105 = io_in_a_bits_opcode == 3'h7;
	wire _T_159 = io_in_a_bits_param != 3'h0;
	wire _T_172 = io_in_a_bits_opcode == 3'h4;
	wire _T_189 = io_in_a_bits_size <= 3'h6;
	wire _T_197 = _T_189 & _T_60;
	wire _T_208 = io_in_a_bits_param == 3'h0;
	wire _T_212 = io_in_a_bits_mask == mask;
	wire _T_220 = io_in_a_bits_opcode == 3'h0;
	wire _T_244 = source_ok & _T_197;
	wire _T_262 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_300 = ~mask;
	wire [3:0] _T_301 = io_in_a_bits_mask & _T_300;
	wire _T_302 = _T_301 == 4'h0;
	wire _T_306 = io_in_a_bits_opcode == 3'h2;
	wire _T_337 = io_in_a_bits_param <= 3'h4;
	wire _T_345 = io_in_a_bits_opcode == 3'h3;
	wire _T_376 = io_in_a_bits_param <= 3'h3;
	wire _T_384 = io_in_a_bits_opcode == 3'h5;
	wire _T_415 = io_in_a_bits_param <= 3'h1;
	wire _T_427 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_431 = io_in_d_bits_opcode == 3'h6;
	wire _T_435 = io_in_d_bits_size >= 3'h2;
	wire _T_439 = io_in_d_bits_param == 2'h0;
	wire _T_443 = ~io_in_d_bits_corrupt;
	wire _T_447 = ~io_in_d_bits_denied;
	wire _T_451 = io_in_d_bits_opcode == 3'h4;
	wire _T_462 = io_in_d_bits_param <= 2'h2;
	wire _T_466 = io_in_d_bits_param != 2'h2;
	wire _T_479 = io_in_d_bits_opcode == 3'h5;
	wire _T_499 = _T_447 | io_in_d_bits_corrupt;
	wire _T_508 = io_in_d_bits_opcode == 3'h0;
	wire _T_525 = io_in_d_bits_opcode == 3'h1;
	wire _T_543 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [3:0] a_first_counter;
	wire [3:0] a_first_counter1 = a_first_counter - 4'h1;
	wire a_first = a_first_counter == 4'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [20:0] address;
	wire _T_573 = io_in_a_valid & ~a_first;
	wire _T_574 = io_in_a_bits_opcode == opcode;
	wire _T_578 = io_in_a_bits_param == param;
	wire _T_582 = io_in_a_bits_size == size;
	wire _T_586 = io_in_a_bits_source == source;
	wire _T_590 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [3:0] d_first_counter;
	wire [3:0] d_first_counter1 = d_first_counter - 4'h1;
	wire d_first = d_first_counter == 4'h0;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_597 = io_in_d_valid & ~d_first;
	wire _T_598 = io_in_d_bits_opcode == opcode_1;
	wire _T_602 = io_in_d_bits_param == param_1;
	wire _T_606 = io_in_d_bits_size == size_1;
	wire _T_610 = io_in_d_bits_source == source_1;
	wire _T_614 = io_in_d_bits_sink == sink;
	wire _T_618 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [3:0] a_first_counter_1;
	wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1;
	wire a_first_1 = a_first_counter_1 == 4'h0;
	reg [3:0] d_first_counter_1;
	wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1;
	wire d_first_1 = d_first_counter_1 == 4'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_624 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire [7:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire _T_627 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_629 = inflight >> io_in_a_bits_source;
	wire _T_631 = ~_T_629[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_635 = io_in_d_valid & d_first_1;
	wire _T_637 = ~_T_431;
	wire _T_638 = (io_in_d_valid & d_first_1) & ~_T_431;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [7:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_431 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_637 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_637 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_624 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_648 = inflight >> io_in_d_bits_source;
	wire _T_650 = _T_648[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_655 = io_in_d_bits_opcode == _GEN_40;
	wire _T_656 = (io_in_d_bits_opcode == _GEN_32) | _T_655;
	wire _T_660 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_667 = io_in_d_bits_opcode == _GEN_56;
	wire _T_668 = (io_in_d_bits_opcode == _GEN_48) | _T_667;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_672 = _GEN_82 == a_size_lookup;
	wire _T_682 = (((_T_635 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_637;
	wire _T_684 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set_wo_ready = _GEN_15[4:0];
	wire [4:0] d_clr_wo_ready = _GEN_21[4:0];
	wire _T_691 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_700 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [3:0] d_first_counter_2;
	wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1;
	wire d_first_2 = d_first_counter_2 == 4'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_726 = (io_in_d_valid & d_first_2) & _T_431;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_431 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_431 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_734 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_744 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_769 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 4'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 4'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 4'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 4'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 4'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 4'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 4'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 4'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 4'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 4'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLFragmenter_7 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [20:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire [7:0] auto_out_a_bits_source;
	output wire [20:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [1:0] auto_out_d_bits_size;
	input [7:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [20:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire repeater_clock;
	wire repeater_reset;
	wire repeater_io_repeat;
	wire repeater_io_full;
	wire repeater_io_enq_ready;
	wire repeater_io_enq_valid;
	wire [2:0] repeater_io_enq_bits_opcode;
	wire [2:0] repeater_io_enq_bits_param;
	wire [2:0] repeater_io_enq_bits_size;
	wire [2:0] repeater_io_enq_bits_source;
	wire [20:0] repeater_io_enq_bits_address;
	wire [3:0] repeater_io_enq_bits_mask;
	wire repeater_io_enq_bits_corrupt;
	wire repeater_io_deq_ready;
	wire repeater_io_deq_valid;
	wire [2:0] repeater_io_deq_bits_opcode;
	wire [2:0] repeater_io_deq_bits_param;
	wire [2:0] repeater_io_deq_bits_size;
	wire [2:0] repeater_io_deq_bits_source;
	wire [20:0] repeater_io_deq_bits_address;
	wire [3:0] repeater_io_deq_bits_mask;
	wire repeater_io_deq_bits_corrupt;
	reg [3:0] acknum;
	reg [2:0] dOrig;
	reg dToggle;
	wire [3:0] dFragnum = auto_out_d_bits_source[3:0];
	wire dFirst = acknum == 4'h0;
	wire dLast = dFragnum == 4'h0;
	wire [3:0] _dsizeOH_T = 4'h1 << auto_out_d_bits_size;
	wire [2:0] dsizeOH = _dsizeOH_T[2:0];
	wire [4:0] _dsizeOH1_T_1 = 5'h03 << auto_out_d_bits_size;
	wire [1:0] dsizeOH1 = ~_dsizeOH1_T_1[1:0];
	wire dHasData = auto_out_d_bits_opcode[0];
	wire _T_5 = ~reset;
	wire ack_decrement = dHasData | dsizeOH[2];
	wire [5:0] _dFirst_size_T = {dFragnum, 2'h0};
	wire [5:0] _GEN_7 = {4'd0, dsizeOH1};
	wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7;
	wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0};
	wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h01;
	wire [6:0] _dFirst_size_T_4 = {1'h0, _dFirst_size_T_1};
	wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4;
	wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5;
	wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4];
	wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0];
	wire _dFirst_size_T_7 = |dFirst_size_hi;
	wire [3:0] _GEN_8 = {1'd0, dFirst_size_hi};
	wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo;
	wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2];
	wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0];
	wire _dFirst_size_T_9 = |dFirst_size_hi_1;
	wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1;
	wire [2:0] dFirst_size = {_dFirst_size_T_7, _dFirst_size_T_9, _dFirst_size_T_10[1]};
	wire drop = ~dHasData & ~dLast;
	wire bundleOut_0_d_ready = auto_in_d_ready | drop;
	wire _T_7 = bundleOut_0_d_ready & auto_out_d_valid;
	wire [3:0] _GEN_9 = {3'd0, ack_decrement};
	wire [3:0] _acknum_T_1 = acknum - _GEN_9;
	wire [2:0] aFrag = (repeater_io_deq_bits_size > 3'h2 ? 3'h2 : repeater_io_deq_bits_size);
	wire [12:0] _aOrigOH1_T_1 = 13'h003f << repeater_io_deq_bits_size;
	wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0];
	wire [8:0] _aFragOH1_T_1 = 9'h003 << aFrag;
	wire [1:0] aFragOH1 = ~_aFragOH1_T_1[1:0];
	wire aHasData = ~repeater_io_deq_bits_opcode[2];
	reg [3:0] gennum;
	wire aFirst = gennum == 4'h0;
	wire [3:0] _old_gennum1_T_2 = gennum - 4'h1;
	wire [3:0] old_gennum1 = (aFirst ? aOrigOH1[5:2] : _old_gennum1_T_2);
	wire [3:0] _new_gennum_T = ~old_gennum1;
	wire [3:0] new_gennum = ~_new_gennum_T;
	reg aToggle_r;
	wire _GEN_5 = (aFirst ? dToggle : aToggle_r);
	wire aToggle = ~_GEN_5;
	wire bundleOut_0_a_valid = repeater_io_deq_valid;
	wire _T_8 = auto_out_a_ready & bundleOut_0_a_valid;
	wire _repeater_io_repeat_T = ~aHasData;
	wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 2'h0};
	wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1;
	wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1;
	wire [5:0] _GEN_10 = {4'd0, aFragOH1};
	wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10;
	wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h03;
	wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4;
	wire [20:0] _GEN_11 = {15'd0, _bundleOut_0_a_bits_address_T_5};
	wire [3:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source, aToggle};
	wire _T_9 = ~repeater_io_full;
	TLMonitor_30 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Repeater_7 repeater(
		.clock(repeater_clock),
		.reset(repeater_reset),
		.io_repeat(repeater_io_repeat),
		.io_full(repeater_io_full),
		.io_enq_ready(repeater_io_enq_ready),
		.io_enq_valid(repeater_io_enq_valid),
		.io_enq_bits_opcode(repeater_io_enq_bits_opcode),
		.io_enq_bits_param(repeater_io_enq_bits_param),
		.io_enq_bits_size(repeater_io_enq_bits_size),
		.io_enq_bits_source(repeater_io_enq_bits_source),
		.io_enq_bits_address(repeater_io_enq_bits_address),
		.io_enq_bits_mask(repeater_io_enq_bits_mask),
		.io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
		.io_deq_ready(repeater_io_deq_ready),
		.io_deq_valid(repeater_io_deq_valid),
		.io_deq_bits_opcode(repeater_io_deq_bits_opcode),
		.io_deq_bits_param(repeater_io_deq_bits_param),
		.io_deq_bits_size(repeater_io_deq_bits_size),
		.io_deq_bits_source(repeater_io_deq_bits_source),
		.io_deq_bits_address(repeater_io_deq_bits_address),
		.io_deq_bits_mask(repeater_io_deq_bits_mask),
		.io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = repeater_io_enq_ready;
	assign auto_in_d_valid = auto_out_d_valid & ~drop;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign auto_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = repeater_io_deq_valid;
	assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode;
	assign auto_out_a_bits_param = repeater_io_deq_bits_param;
	assign auto_out_a_bits_size = aFrag[1:0];
	assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi, new_gennum};
	assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11;
	assign auto_out_a_bits_mask = (repeater_io_full ? 4'hf : auto_in_a_bits_mask);
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready | drop;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = repeater_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid & ~drop;
	assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_io_in_d_bits_param = auto_out_d_bits_param;
	assign monitor_io_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign monitor_io_in_d_bits_source = auto_out_d_bits_source[7:5];
	assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink;
	assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied;
	assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign repeater_clock = clock;
	assign repeater_reset = reset;
	assign repeater_io_repeat = ~aHasData & (new_gennum != 4'h0);
	assign repeater_io_enq_valid = auto_in_a_valid;
	assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign repeater_io_enq_bits_param = auto_in_a_bits_param;
	assign repeater_io_enq_bits_size = auto_in_a_bits_size;
	assign repeater_io_enq_bits_source = auto_in_a_bits_source;
	assign repeater_io_enq_bits_address = auto_in_a_bits_address;
	assign repeater_io_enq_bits_mask = auto_in_a_bits_mask;
	assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign repeater_io_deq_ready = auto_out_a_ready;
	always @(posedge clock) begin
		if (reset)
			acknum <= 4'h0;
		else if (_T_7)
			if (dFirst)
				acknum <= dFragnum;
			else
				acknum <= _acknum_T_1;
		if (_T_7)
			if (dFirst)
				dOrig <= dFirst_size;
		if (reset)
			dToggle <= 1'h0;
		else if (_T_7)
			if (dFirst)
				dToggle <= auto_out_d_bits_source[4];
		if (reset)
			gennum <= 4'h0;
		else if (_T_8)
			gennum <= new_gennum;
		if (aFirst)
			aToggle_r <= dToggle;
	end
endmodule
module TLInterconnectCoupler_17 (
	clock,
	reset,
	auto_buffer_in_a_ready,
	auto_buffer_in_a_valid,
	auto_buffer_in_a_bits_opcode,
	auto_buffer_in_a_bits_param,
	auto_buffer_in_a_bits_size,
	auto_buffer_in_a_bits_source,
	auto_buffer_in_a_bits_address,
	auto_buffer_in_a_bits_mask,
	auto_buffer_in_a_bits_data,
	auto_buffer_in_a_bits_corrupt,
	auto_buffer_in_d_ready,
	auto_buffer_in_d_valid,
	auto_buffer_in_d_bits_opcode,
	auto_buffer_in_d_bits_param,
	auto_buffer_in_d_bits_size,
	auto_buffer_in_d_bits_source,
	auto_buffer_in_d_bits_sink,
	auto_buffer_in_d_bits_denied,
	auto_buffer_in_d_bits_data,
	auto_buffer_in_d_bits_corrupt,
	auto_buffer_out_a_ready,
	auto_buffer_out_a_valid,
	auto_buffer_out_a_bits_opcode,
	auto_buffer_out_a_bits_param,
	auto_buffer_out_a_bits_size,
	auto_buffer_out_a_bits_source,
	auto_buffer_out_a_bits_address,
	auto_buffer_out_a_bits_mask,
	auto_buffer_out_a_bits_data,
	auto_buffer_out_a_bits_corrupt,
	auto_buffer_out_d_ready,
	auto_buffer_out_d_valid,
	auto_buffer_out_d_bits_opcode,
	auto_buffer_out_d_bits_size,
	auto_buffer_out_d_bits_source,
	auto_buffer_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_buffer_in_a_ready;
	input auto_buffer_in_a_valid;
	input [2:0] auto_buffer_in_a_bits_opcode;
	input [2:0] auto_buffer_in_a_bits_param;
	input [2:0] auto_buffer_in_a_bits_size;
	input [2:0] auto_buffer_in_a_bits_source;
	input [20:0] auto_buffer_in_a_bits_address;
	input [3:0] auto_buffer_in_a_bits_mask;
	input [31:0] auto_buffer_in_a_bits_data;
	input auto_buffer_in_a_bits_corrupt;
	input auto_buffer_in_d_ready;
	output wire auto_buffer_in_d_valid;
	output wire [2:0] auto_buffer_in_d_bits_opcode;
	output wire [1:0] auto_buffer_in_d_bits_param;
	output wire [2:0] auto_buffer_in_d_bits_size;
	output wire [2:0] auto_buffer_in_d_bits_source;
	output wire auto_buffer_in_d_bits_sink;
	output wire auto_buffer_in_d_bits_denied;
	output wire [31:0] auto_buffer_in_d_bits_data;
	output wire auto_buffer_in_d_bits_corrupt;
	input auto_buffer_out_a_ready;
	output wire auto_buffer_out_a_valid;
	output wire [2:0] auto_buffer_out_a_bits_opcode;
	output wire [2:0] auto_buffer_out_a_bits_param;
	output wire [1:0] auto_buffer_out_a_bits_size;
	output wire [7:0] auto_buffer_out_a_bits_source;
	output wire [20:0] auto_buffer_out_a_bits_address;
	output wire [3:0] auto_buffer_out_a_bits_mask;
	output wire [31:0] auto_buffer_out_a_bits_data;
	output wire auto_buffer_out_a_bits_corrupt;
	output wire auto_buffer_out_d_ready;
	input auto_buffer_out_d_valid;
	input [2:0] auto_buffer_out_d_bits_opcode;
	input [1:0] auto_buffer_out_d_bits_size;
	input [7:0] auto_buffer_out_d_bits_source;
	input [31:0] auto_buffer_out_d_bits_data;
	wire buffer_clock;
	wire buffer_reset;
	wire buffer_auto_in_a_ready;
	wire buffer_auto_in_a_valid;
	wire [2:0] buffer_auto_in_a_bits_opcode;
	wire [2:0] buffer_auto_in_a_bits_param;
	wire [1:0] buffer_auto_in_a_bits_size;
	wire [7:0] buffer_auto_in_a_bits_source;
	wire [20:0] buffer_auto_in_a_bits_address;
	wire [3:0] buffer_auto_in_a_bits_mask;
	wire [31:0] buffer_auto_in_a_bits_data;
	wire buffer_auto_in_a_bits_corrupt;
	wire buffer_auto_in_d_ready;
	wire buffer_auto_in_d_valid;
	wire [2:0] buffer_auto_in_d_bits_opcode;
	wire [1:0] buffer_auto_in_d_bits_param;
	wire [1:0] buffer_auto_in_d_bits_size;
	wire [7:0] buffer_auto_in_d_bits_source;
	wire buffer_auto_in_d_bits_sink;
	wire buffer_auto_in_d_bits_denied;
	wire [31:0] buffer_auto_in_d_bits_data;
	wire buffer_auto_in_d_bits_corrupt;
	wire buffer_auto_out_a_ready;
	wire buffer_auto_out_a_valid;
	wire [2:0] buffer_auto_out_a_bits_opcode;
	wire [2:0] buffer_auto_out_a_bits_param;
	wire [1:0] buffer_auto_out_a_bits_size;
	wire [7:0] buffer_auto_out_a_bits_source;
	wire [20:0] buffer_auto_out_a_bits_address;
	wire [3:0] buffer_auto_out_a_bits_mask;
	wire [31:0] buffer_auto_out_a_bits_data;
	wire buffer_auto_out_a_bits_corrupt;
	wire buffer_auto_out_d_ready;
	wire buffer_auto_out_d_valid;
	wire [2:0] buffer_auto_out_d_bits_opcode;
	wire [1:0] buffer_auto_out_d_bits_size;
	wire [7:0] buffer_auto_out_d_bits_source;
	wire [31:0] buffer_auto_out_d_bits_data;
	wire fragmenter_clock;
	wire fragmenter_reset;
	wire fragmenter_auto_in_a_ready;
	wire fragmenter_auto_in_a_valid;
	wire [2:0] fragmenter_auto_in_a_bits_opcode;
	wire [2:0] fragmenter_auto_in_a_bits_param;
	wire [2:0] fragmenter_auto_in_a_bits_size;
	wire [2:0] fragmenter_auto_in_a_bits_source;
	wire [20:0] fragmenter_auto_in_a_bits_address;
	wire [3:0] fragmenter_auto_in_a_bits_mask;
	wire [31:0] fragmenter_auto_in_a_bits_data;
	wire fragmenter_auto_in_a_bits_corrupt;
	wire fragmenter_auto_in_d_ready;
	wire fragmenter_auto_in_d_valid;
	wire [2:0] fragmenter_auto_in_d_bits_opcode;
	wire [1:0] fragmenter_auto_in_d_bits_param;
	wire [2:0] fragmenter_auto_in_d_bits_size;
	wire [2:0] fragmenter_auto_in_d_bits_source;
	wire fragmenter_auto_in_d_bits_sink;
	wire fragmenter_auto_in_d_bits_denied;
	wire [31:0] fragmenter_auto_in_d_bits_data;
	wire fragmenter_auto_in_d_bits_corrupt;
	wire fragmenter_auto_out_a_ready;
	wire fragmenter_auto_out_a_valid;
	wire [2:0] fragmenter_auto_out_a_bits_opcode;
	wire [2:0] fragmenter_auto_out_a_bits_param;
	wire [1:0] fragmenter_auto_out_a_bits_size;
	wire [7:0] fragmenter_auto_out_a_bits_source;
	wire [20:0] fragmenter_auto_out_a_bits_address;
	wire [3:0] fragmenter_auto_out_a_bits_mask;
	wire [31:0] fragmenter_auto_out_a_bits_data;
	wire fragmenter_auto_out_a_bits_corrupt;
	wire fragmenter_auto_out_d_ready;
	wire fragmenter_auto_out_d_valid;
	wire [2:0] fragmenter_auto_out_d_bits_opcode;
	wire [1:0] fragmenter_auto_out_d_bits_param;
	wire [1:0] fragmenter_auto_out_d_bits_size;
	wire [7:0] fragmenter_auto_out_d_bits_source;
	wire fragmenter_auto_out_d_bits_sink;
	wire fragmenter_auto_out_d_bits_denied;
	wire [31:0] fragmenter_auto_out_d_bits_data;
	wire fragmenter_auto_out_d_bits_corrupt;
	wire buffer_1_auto_in_a_ready;
	wire buffer_1_auto_in_a_valid;
	wire [2:0] buffer_1_auto_in_a_bits_opcode;
	wire [2:0] buffer_1_auto_in_a_bits_param;
	wire [2:0] buffer_1_auto_in_a_bits_size;
	wire [2:0] buffer_1_auto_in_a_bits_source;
	wire [20:0] buffer_1_auto_in_a_bits_address;
	wire [3:0] buffer_1_auto_in_a_bits_mask;
	wire [31:0] buffer_1_auto_in_a_bits_data;
	wire buffer_1_auto_in_a_bits_corrupt;
	wire buffer_1_auto_in_d_ready;
	wire buffer_1_auto_in_d_valid;
	wire [2:0] buffer_1_auto_in_d_bits_opcode;
	wire [1:0] buffer_1_auto_in_d_bits_param;
	wire [2:0] buffer_1_auto_in_d_bits_size;
	wire [2:0] buffer_1_auto_in_d_bits_source;
	wire buffer_1_auto_in_d_bits_sink;
	wire buffer_1_auto_in_d_bits_denied;
	wire [31:0] buffer_1_auto_in_d_bits_data;
	wire buffer_1_auto_in_d_bits_corrupt;
	wire buffer_1_auto_out_a_ready;
	wire buffer_1_auto_out_a_valid;
	wire [2:0] buffer_1_auto_out_a_bits_opcode;
	wire [2:0] buffer_1_auto_out_a_bits_param;
	wire [2:0] buffer_1_auto_out_a_bits_size;
	wire [2:0] buffer_1_auto_out_a_bits_source;
	wire [20:0] buffer_1_auto_out_a_bits_address;
	wire [3:0] buffer_1_auto_out_a_bits_mask;
	wire [31:0] buffer_1_auto_out_a_bits_data;
	wire buffer_1_auto_out_a_bits_corrupt;
	wire buffer_1_auto_out_d_ready;
	wire buffer_1_auto_out_d_valid;
	wire [2:0] buffer_1_auto_out_d_bits_opcode;
	wire [1:0] buffer_1_auto_out_d_bits_param;
	wire [2:0] buffer_1_auto_out_d_bits_size;
	wire [2:0] buffer_1_auto_out_d_bits_source;
	wire buffer_1_auto_out_d_bits_sink;
	wire buffer_1_auto_out_d_bits_denied;
	wire [31:0] buffer_1_auto_out_d_bits_data;
	wire buffer_1_auto_out_d_bits_corrupt;
	TLBuffer_11 buffer(
		.clock(buffer_clock),
		.reset(buffer_reset),
		.auto_in_a_ready(buffer_auto_in_a_ready),
		.auto_in_a_valid(buffer_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_auto_in_d_ready),
		.auto_in_d_valid(buffer_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_auto_out_a_ready),
		.auto_out_a_valid(buffer_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_auto_out_d_ready),
		.auto_out_d_valid(buffer_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(buffer_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_auto_out_d_bits_source),
		.auto_out_d_bits_data(buffer_auto_out_d_bits_data)
	);
	TLFragmenter_7 fragmenter(
		.clock(fragmenter_clock),
		.reset(fragmenter_reset),
		.auto_in_a_ready(fragmenter_auto_in_a_ready),
		.auto_in_a_valid(fragmenter_auto_in_a_valid),
		.auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
		.auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
		.auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
		.auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
		.auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
		.auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
		.auto_in_d_ready(fragmenter_auto_in_d_ready),
		.auto_in_d_valid(fragmenter_auto_in_d_valid),
		.auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(fragmenter_auto_in_d_bits_param),
		.auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
		.auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
		.auto_in_d_bits_sink(fragmenter_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(fragmenter_auto_in_d_bits_denied),
		.auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(fragmenter_auto_in_d_bits_corrupt),
		.auto_out_a_ready(fragmenter_auto_out_a_ready),
		.auto_out_a_valid(fragmenter_auto_out_a_valid),
		.auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
		.auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
		.auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
		.auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
		.auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
		.auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
		.auto_out_d_ready(fragmenter_auto_out_d_ready),
		.auto_out_d_valid(fragmenter_auto_out_d_valid),
		.auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(fragmenter_auto_out_d_bits_param),
		.auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
		.auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
		.auto_out_d_bits_sink(fragmenter_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(fragmenter_auto_out_d_bits_denied),
		.auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(fragmenter_auto_out_d_bits_corrupt)
	);
	TLBuffer_10 buffer_1(
		.auto_in_a_ready(buffer_1_auto_in_a_ready),
		.auto_in_a_valid(buffer_1_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_1_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_1_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_1_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_1_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_1_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_1_auto_in_d_ready),
		.auto_in_d_valid(buffer_1_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_1_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_1_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_1_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_1_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_1_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_1_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_1_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_1_auto_out_a_ready),
		.auto_out_a_valid(buffer_1_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_1_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_1_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_1_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_1_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_1_auto_out_d_ready),
		.auto_out_d_valid(buffer_1_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(buffer_1_auto_out_d_bits_param),
		.auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
		.auto_out_d_bits_sink(buffer_1_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
		.auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt)
	);
	assign auto_buffer_in_a_ready = buffer_1_auto_in_a_ready;
	assign auto_buffer_in_d_valid = buffer_1_auto_in_d_valid;
	assign auto_buffer_in_d_bits_opcode = buffer_1_auto_in_d_bits_opcode;
	assign auto_buffer_in_d_bits_param = buffer_1_auto_in_d_bits_param;
	assign auto_buffer_in_d_bits_size = buffer_1_auto_in_d_bits_size;
	assign auto_buffer_in_d_bits_source = buffer_1_auto_in_d_bits_source;
	assign auto_buffer_in_d_bits_sink = buffer_1_auto_in_d_bits_sink;
	assign auto_buffer_in_d_bits_denied = buffer_1_auto_in_d_bits_denied;
	assign auto_buffer_in_d_bits_data = buffer_1_auto_in_d_bits_data;
	assign auto_buffer_in_d_bits_corrupt = buffer_1_auto_in_d_bits_corrupt;
	assign auto_buffer_out_a_valid = buffer_auto_out_a_valid;
	assign auto_buffer_out_a_bits_opcode = buffer_auto_out_a_bits_opcode;
	assign auto_buffer_out_a_bits_param = buffer_auto_out_a_bits_param;
	assign auto_buffer_out_a_bits_size = buffer_auto_out_a_bits_size;
	assign auto_buffer_out_a_bits_source = buffer_auto_out_a_bits_source;
	assign auto_buffer_out_a_bits_address = buffer_auto_out_a_bits_address;
	assign auto_buffer_out_a_bits_mask = buffer_auto_out_a_bits_mask;
	assign auto_buffer_out_a_bits_data = buffer_auto_out_a_bits_data;
	assign auto_buffer_out_a_bits_corrupt = buffer_auto_out_a_bits_corrupt;
	assign auto_buffer_out_d_ready = buffer_auto_out_d_ready;
	assign buffer_clock = clock;
	assign buffer_reset = reset;
	assign buffer_auto_in_a_valid = fragmenter_auto_out_a_valid;
	assign buffer_auto_in_a_bits_opcode = fragmenter_auto_out_a_bits_opcode;
	assign buffer_auto_in_a_bits_param = fragmenter_auto_out_a_bits_param;
	assign buffer_auto_in_a_bits_size = fragmenter_auto_out_a_bits_size;
	assign buffer_auto_in_a_bits_source = fragmenter_auto_out_a_bits_source;
	assign buffer_auto_in_a_bits_address = fragmenter_auto_out_a_bits_address;
	assign buffer_auto_in_a_bits_mask = fragmenter_auto_out_a_bits_mask;
	assign buffer_auto_in_a_bits_data = fragmenter_auto_out_a_bits_data;
	assign buffer_auto_in_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt;
	assign buffer_auto_in_d_ready = fragmenter_auto_out_d_ready;
	assign buffer_auto_out_a_ready = auto_buffer_out_a_ready;
	assign buffer_auto_out_d_valid = auto_buffer_out_d_valid;
	assign buffer_auto_out_d_bits_opcode = auto_buffer_out_d_bits_opcode;
	assign buffer_auto_out_d_bits_size = auto_buffer_out_d_bits_size;
	assign buffer_auto_out_d_bits_source = auto_buffer_out_d_bits_source;
	assign buffer_auto_out_d_bits_data = auto_buffer_out_d_bits_data;
	assign fragmenter_clock = clock;
	assign fragmenter_reset = reset;
	assign fragmenter_auto_in_a_valid = buffer_1_auto_out_a_valid;
	assign fragmenter_auto_in_a_bits_opcode = buffer_1_auto_out_a_bits_opcode;
	assign fragmenter_auto_in_a_bits_param = buffer_1_auto_out_a_bits_param;
	assign fragmenter_auto_in_a_bits_size = buffer_1_auto_out_a_bits_size;
	assign fragmenter_auto_in_a_bits_source = buffer_1_auto_out_a_bits_source;
	assign fragmenter_auto_in_a_bits_address = buffer_1_auto_out_a_bits_address;
	assign fragmenter_auto_in_a_bits_mask = buffer_1_auto_out_a_bits_mask;
	assign fragmenter_auto_in_a_bits_data = buffer_1_auto_out_a_bits_data;
	assign fragmenter_auto_in_a_bits_corrupt = buffer_1_auto_out_a_bits_corrupt;
	assign fragmenter_auto_in_d_ready = buffer_1_auto_out_d_ready;
	assign fragmenter_auto_out_a_ready = buffer_auto_in_a_ready;
	assign fragmenter_auto_out_d_valid = buffer_auto_in_d_valid;
	assign fragmenter_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode;
	assign fragmenter_auto_out_d_bits_param = buffer_auto_in_d_bits_param;
	assign fragmenter_auto_out_d_bits_size = buffer_auto_in_d_bits_size;
	assign fragmenter_auto_out_d_bits_source = buffer_auto_in_d_bits_source;
	assign fragmenter_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink;
	assign fragmenter_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied;
	assign fragmenter_auto_out_d_bits_data = buffer_auto_in_d_bits_data;
	assign fragmenter_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt;
	assign buffer_1_auto_in_a_valid = auto_buffer_in_a_valid;
	assign buffer_1_auto_in_a_bits_opcode = auto_buffer_in_a_bits_opcode;
	assign buffer_1_auto_in_a_bits_param = auto_buffer_in_a_bits_param;
	assign buffer_1_auto_in_a_bits_size = auto_buffer_in_a_bits_size;
	assign buffer_1_auto_in_a_bits_source = auto_buffer_in_a_bits_source;
	assign buffer_1_auto_in_a_bits_address = auto_buffer_in_a_bits_address;
	assign buffer_1_auto_in_a_bits_mask = auto_buffer_in_a_bits_mask;
	assign buffer_1_auto_in_a_bits_data = auto_buffer_in_a_bits_data;
	assign buffer_1_auto_in_a_bits_corrupt = auto_buffer_in_a_bits_corrupt;
	assign buffer_1_auto_in_d_ready = auto_buffer_in_d_ready;
	assign buffer_1_auto_out_a_ready = fragmenter_auto_in_a_ready;
	assign buffer_1_auto_out_d_valid = fragmenter_auto_in_d_valid;
	assign buffer_1_auto_out_d_bits_opcode = fragmenter_auto_in_d_bits_opcode;
	assign buffer_1_auto_out_d_bits_param = fragmenter_auto_in_d_bits_param;
	assign buffer_1_auto_out_d_bits_size = fragmenter_auto_in_d_bits_size;
	assign buffer_1_auto_out_d_bits_source = fragmenter_auto_in_d_bits_source;
	assign buffer_1_auto_out_d_bits_sink = fragmenter_auto_in_d_bits_sink;
	assign buffer_1_auto_out_d_bits_denied = fragmenter_auto_in_d_bits_denied;
	assign buffer_1_auto_out_d_bits_data = fragmenter_auto_in_d_bits_data;
	assign buffer_1_auto_out_d_bits_corrupt = fragmenter_auto_in_d_bits_corrupt;
endmodule
module PeripheryBus_1 (
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_ready,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_valid,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_opcode,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_param,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_size,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_source,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_address,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_mask,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_data,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_corrupt,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_ready,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_valid,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_opcode,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_size,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_source,
	auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_data,
	auto_coupler_to_slave_named_clockgater_buffer_out_a_ready,
	auto_coupler_to_slave_named_clockgater_buffer_out_a_valid,
	auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_opcode,
	auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_param,
	auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_size,
	auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_source,
	auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_address,
	auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_mask,
	auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_data,
	auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_corrupt,
	auto_coupler_to_slave_named_clockgater_buffer_out_d_ready,
	auto_coupler_to_slave_named_clockgater_buffer_out_d_valid,
	auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_opcode,
	auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_size,
	auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_source,
	auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_data,
	auto_coupler_to_bootrom_fragmenter_out_a_ready,
	auto_coupler_to_bootrom_fragmenter_out_a_valid,
	auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode,
	auto_coupler_to_bootrom_fragmenter_out_a_bits_param,
	auto_coupler_to_bootrom_fragmenter_out_a_bits_size,
	auto_coupler_to_bootrom_fragmenter_out_a_bits_source,
	auto_coupler_to_bootrom_fragmenter_out_a_bits_address,
	auto_coupler_to_bootrom_fragmenter_out_a_bits_mask,
	auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt,
	auto_coupler_to_bootrom_fragmenter_out_d_ready,
	auto_coupler_to_bootrom_fragmenter_out_d_valid,
	auto_coupler_to_bootrom_fragmenter_out_d_bits_size,
	auto_coupler_to_bootrom_fragmenter_out_d_bits_source,
	auto_coupler_to_bootrom_fragmenter_out_d_bits_data,
	auto_coupler_to_tile_tl_slave_clock_xing_out_a_ready,
	auto_coupler_to_tile_tl_slave_clock_xing_out_a_valid,
	auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_opcode,
	auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_param,
	auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_size,
	auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_source,
	auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_address,
	auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_mask,
	auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_data,
	auto_coupler_to_tile_tl_slave_clock_xing_out_d_ready,
	auto_coupler_to_tile_tl_slave_clock_xing_out_d_valid,
	auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_opcode,
	auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_param,
	auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_size,
	auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_source,
	auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_sink,
	auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_denied,
	auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_data,
	auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_corrupt,
	auto_coupler_to_debug_fragmenter_out_a_ready,
	auto_coupler_to_debug_fragmenter_out_a_valid,
	auto_coupler_to_debug_fragmenter_out_a_bits_opcode,
	auto_coupler_to_debug_fragmenter_out_a_bits_param,
	auto_coupler_to_debug_fragmenter_out_a_bits_size,
	auto_coupler_to_debug_fragmenter_out_a_bits_source,
	auto_coupler_to_debug_fragmenter_out_a_bits_address,
	auto_coupler_to_debug_fragmenter_out_a_bits_mask,
	auto_coupler_to_debug_fragmenter_out_a_bits_data,
	auto_coupler_to_debug_fragmenter_out_a_bits_corrupt,
	auto_coupler_to_debug_fragmenter_out_d_ready,
	auto_coupler_to_debug_fragmenter_out_d_valid,
	auto_coupler_to_debug_fragmenter_out_d_bits_opcode,
	auto_coupler_to_debug_fragmenter_out_d_bits_size,
	auto_coupler_to_debug_fragmenter_out_d_bits_source,
	auto_coupler_to_debug_fragmenter_out_d_bits_data,
	auto_coupler_to_clint_fragmenter_out_a_ready,
	auto_coupler_to_clint_fragmenter_out_a_valid,
	auto_coupler_to_clint_fragmenter_out_a_bits_opcode,
	auto_coupler_to_clint_fragmenter_out_a_bits_param,
	auto_coupler_to_clint_fragmenter_out_a_bits_size,
	auto_coupler_to_clint_fragmenter_out_a_bits_source,
	auto_coupler_to_clint_fragmenter_out_a_bits_address,
	auto_coupler_to_clint_fragmenter_out_a_bits_mask,
	auto_coupler_to_clint_fragmenter_out_a_bits_data,
	auto_coupler_to_clint_fragmenter_out_a_bits_corrupt,
	auto_coupler_to_clint_fragmenter_out_d_ready,
	auto_coupler_to_clint_fragmenter_out_d_valid,
	auto_coupler_to_clint_fragmenter_out_d_bits_opcode,
	auto_coupler_to_clint_fragmenter_out_d_bits_size,
	auto_coupler_to_clint_fragmenter_out_d_bits_source,
	auto_coupler_to_clint_fragmenter_out_d_bits_data,
	auto_coupler_to_plic_fragmenter_out_a_ready,
	auto_coupler_to_plic_fragmenter_out_a_valid,
	auto_coupler_to_plic_fragmenter_out_a_bits_opcode,
	auto_coupler_to_plic_fragmenter_out_a_bits_param,
	auto_coupler_to_plic_fragmenter_out_a_bits_size,
	auto_coupler_to_plic_fragmenter_out_a_bits_source,
	auto_coupler_to_plic_fragmenter_out_a_bits_address,
	auto_coupler_to_plic_fragmenter_out_a_bits_mask,
	auto_coupler_to_plic_fragmenter_out_a_bits_data,
	auto_coupler_to_plic_fragmenter_out_a_bits_corrupt,
	auto_coupler_to_plic_fragmenter_out_d_ready,
	auto_coupler_to_plic_fragmenter_out_d_valid,
	auto_coupler_to_plic_fragmenter_out_d_bits_opcode,
	auto_coupler_to_plic_fragmenter_out_d_bits_size,
	auto_coupler_to_plic_fragmenter_out_d_bits_source,
	auto_coupler_to_plic_fragmenter_out_d_bits_data,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_corrupt,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_param,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_sink,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data,
	auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt,
	auto_fixedClockNode_out_4_clock,
	auto_fixedClockNode_out_4_reset,
	auto_fixedClockNode_out_3_clock,
	auto_fixedClockNode_out_3_reset,
	auto_fixedClockNode_out_2_clock,
	auto_fixedClockNode_out_2_reset,
	auto_fixedClockNode_out_0_clock,
	auto_fixedClockNode_out_0_reset,
	auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock,
	auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset,
	auto_bus_xing_in_a_ready,
	auto_bus_xing_in_a_valid,
	auto_bus_xing_in_a_bits_opcode,
	auto_bus_xing_in_a_bits_param,
	auto_bus_xing_in_a_bits_size,
	auto_bus_xing_in_a_bits_source,
	auto_bus_xing_in_a_bits_address,
	auto_bus_xing_in_a_bits_mask,
	auto_bus_xing_in_a_bits_data,
	auto_bus_xing_in_a_bits_corrupt,
	auto_bus_xing_in_d_ready,
	auto_bus_xing_in_d_valid,
	auto_bus_xing_in_d_bits_opcode,
	auto_bus_xing_in_d_bits_param,
	auto_bus_xing_in_d_bits_size,
	auto_bus_xing_in_d_bits_source,
	auto_bus_xing_in_d_bits_sink,
	auto_bus_xing_in_d_bits_denied,
	auto_bus_xing_in_d_bits_data,
	auto_bus_xing_in_d_bits_corrupt,
	custom_boot,
	clock,
	reset
);
	input auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_ready;
	output wire auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_valid;
	output wire [2:0] auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_opcode;
	output wire [2:0] auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_param;
	output wire [1:0] auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_size;
	output wire [7:0] auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_source;
	output wire [20:0] auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_address;
	output wire [3:0] auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_mask;
	output wire [31:0] auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_data;
	output wire auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_corrupt;
	output wire auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_ready;
	input auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_valid;
	input [2:0] auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_opcode;
	input [1:0] auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_size;
	input [7:0] auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_source;
	input [31:0] auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_data;
	input auto_coupler_to_slave_named_clockgater_buffer_out_a_ready;
	output wire auto_coupler_to_slave_named_clockgater_buffer_out_a_valid;
	output wire [2:0] auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_opcode;
	output wire [2:0] auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_param;
	output wire [1:0] auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_size;
	output wire [7:0] auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_source;
	output wire [20:0] auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_address;
	output wire [3:0] auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_mask;
	output wire [31:0] auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_data;
	output wire auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_corrupt;
	output wire auto_coupler_to_slave_named_clockgater_buffer_out_d_ready;
	input auto_coupler_to_slave_named_clockgater_buffer_out_d_valid;
	input [2:0] auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_opcode;
	input [1:0] auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_size;
	input [7:0] auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_source;
	input [31:0] auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_data;
	input auto_coupler_to_bootrom_fragmenter_out_a_ready;
	output wire auto_coupler_to_bootrom_fragmenter_out_a_valid;
	output wire [2:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode;
	output wire [2:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_param;
	output wire [1:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_size;
	output wire [7:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_source;
	output wire [16:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_address;
	output wire [3:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_mask;
	output wire auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt;
	output wire auto_coupler_to_bootrom_fragmenter_out_d_ready;
	input auto_coupler_to_bootrom_fragmenter_out_d_valid;
	input [1:0] auto_coupler_to_bootrom_fragmenter_out_d_bits_size;
	input [7:0] auto_coupler_to_bootrom_fragmenter_out_d_bits_source;
	input [31:0] auto_coupler_to_bootrom_fragmenter_out_d_bits_data;
	input auto_coupler_to_tile_tl_slave_clock_xing_out_a_ready;
	output wire auto_coupler_to_tile_tl_slave_clock_xing_out_a_valid;
	output wire [2:0] auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_opcode;
	output wire [2:0] auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_param;
	output wire [2:0] auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_size;
	output wire [2:0] auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_source;
	output wire [31:0] auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_address;
	output wire [3:0] auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_mask;
	output wire [31:0] auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_data;
	output wire auto_coupler_to_tile_tl_slave_clock_xing_out_d_ready;
	input auto_coupler_to_tile_tl_slave_clock_xing_out_d_valid;
	input [2:0] auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_opcode;
	input [1:0] auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_param;
	input [2:0] auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_size;
	input [2:0] auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_source;
	input auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_sink;
	input auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_denied;
	input [31:0] auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_data;
	input auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_corrupt;
	input auto_coupler_to_debug_fragmenter_out_a_ready;
	output wire auto_coupler_to_debug_fragmenter_out_a_valid;
	output wire [2:0] auto_coupler_to_debug_fragmenter_out_a_bits_opcode;
	output wire [2:0] auto_coupler_to_debug_fragmenter_out_a_bits_param;
	output wire [1:0] auto_coupler_to_debug_fragmenter_out_a_bits_size;
	output wire [7:0] auto_coupler_to_debug_fragmenter_out_a_bits_source;
	output wire [11:0] auto_coupler_to_debug_fragmenter_out_a_bits_address;
	output wire [3:0] auto_coupler_to_debug_fragmenter_out_a_bits_mask;
	output wire [31:0] auto_coupler_to_debug_fragmenter_out_a_bits_data;
	output wire auto_coupler_to_debug_fragmenter_out_a_bits_corrupt;
	output wire auto_coupler_to_debug_fragmenter_out_d_ready;
	input auto_coupler_to_debug_fragmenter_out_d_valid;
	input [2:0] auto_coupler_to_debug_fragmenter_out_d_bits_opcode;
	input [1:0] auto_coupler_to_debug_fragmenter_out_d_bits_size;
	input [7:0] auto_coupler_to_debug_fragmenter_out_d_bits_source;
	input [31:0] auto_coupler_to_debug_fragmenter_out_d_bits_data;
	input auto_coupler_to_clint_fragmenter_out_a_ready;
	output wire auto_coupler_to_clint_fragmenter_out_a_valid;
	output wire [2:0] auto_coupler_to_clint_fragmenter_out_a_bits_opcode;
	output wire [2:0] auto_coupler_to_clint_fragmenter_out_a_bits_param;
	output wire [1:0] auto_coupler_to_clint_fragmenter_out_a_bits_size;
	output wire [7:0] auto_coupler_to_clint_fragmenter_out_a_bits_source;
	output wire [25:0] auto_coupler_to_clint_fragmenter_out_a_bits_address;
	output wire [3:0] auto_coupler_to_clint_fragmenter_out_a_bits_mask;
	output wire [31:0] auto_coupler_to_clint_fragmenter_out_a_bits_data;
	output wire auto_coupler_to_clint_fragmenter_out_a_bits_corrupt;
	output wire auto_coupler_to_clint_fragmenter_out_d_ready;
	input auto_coupler_to_clint_fragmenter_out_d_valid;
	input [2:0] auto_coupler_to_clint_fragmenter_out_d_bits_opcode;
	input [1:0] auto_coupler_to_clint_fragmenter_out_d_bits_size;
	input [7:0] auto_coupler_to_clint_fragmenter_out_d_bits_source;
	input [31:0] auto_coupler_to_clint_fragmenter_out_d_bits_data;
	input auto_coupler_to_plic_fragmenter_out_a_ready;
	output wire auto_coupler_to_plic_fragmenter_out_a_valid;
	output wire [2:0] auto_coupler_to_plic_fragmenter_out_a_bits_opcode;
	output wire [2:0] auto_coupler_to_plic_fragmenter_out_a_bits_param;
	output wire [1:0] auto_coupler_to_plic_fragmenter_out_a_bits_size;
	output wire [7:0] auto_coupler_to_plic_fragmenter_out_a_bits_source;
	output wire [27:0] auto_coupler_to_plic_fragmenter_out_a_bits_address;
	output wire [3:0] auto_coupler_to_plic_fragmenter_out_a_bits_mask;
	output wire [31:0] auto_coupler_to_plic_fragmenter_out_a_bits_data;
	output wire auto_coupler_to_plic_fragmenter_out_a_bits_corrupt;
	output wire auto_coupler_to_plic_fragmenter_out_d_ready;
	input auto_coupler_to_plic_fragmenter_out_d_valid;
	input [2:0] auto_coupler_to_plic_fragmenter_out_d_bits_opcode;
	input [1:0] auto_coupler_to_plic_fragmenter_out_d_bits_size;
	input [7:0] auto_coupler_to_plic_fragmenter_out_d_bits_source;
	input [31:0] auto_coupler_to_plic_fragmenter_out_d_bits_data;
	input auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready;
	output wire auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid;
	output wire [2:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode;
	output wire [2:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param;
	output wire [2:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size;
	output wire [2:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source;
	output wire [30:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address;
	output wire [3:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask;
	output wire [31:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data;
	output wire auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_corrupt;
	output wire auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready;
	input auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid;
	input [2:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode;
	input [1:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_param;
	input [2:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size;
	input [2:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source;
	input auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_sink;
	input auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied;
	input [31:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data;
	input auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt;
	output wire auto_fixedClockNode_out_4_clock;
	output wire auto_fixedClockNode_out_4_reset;
	output wire auto_fixedClockNode_out_3_clock;
	output wire auto_fixedClockNode_out_3_reset;
	output wire auto_fixedClockNode_out_2_clock;
	output wire auto_fixedClockNode_out_2_reset;
	output wire auto_fixedClockNode_out_0_clock;
	output wire auto_fixedClockNode_out_0_reset;
	input auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock;
	input auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset;
	output wire auto_bus_xing_in_a_ready;
	input auto_bus_xing_in_a_valid;
	input [2:0] auto_bus_xing_in_a_bits_opcode;
	input [2:0] auto_bus_xing_in_a_bits_param;
	input [3:0] auto_bus_xing_in_a_bits_size;
	input [1:0] auto_bus_xing_in_a_bits_source;
	input [31:0] auto_bus_xing_in_a_bits_address;
	input [3:0] auto_bus_xing_in_a_bits_mask;
	input [31:0] auto_bus_xing_in_a_bits_data;
	input auto_bus_xing_in_a_bits_corrupt;
	input auto_bus_xing_in_d_ready;
	output wire auto_bus_xing_in_d_valid;
	output wire [2:0] auto_bus_xing_in_d_bits_opcode;
	output wire [1:0] auto_bus_xing_in_d_bits_param;
	output wire [3:0] auto_bus_xing_in_d_bits_size;
	output wire [1:0] auto_bus_xing_in_d_bits_source;
	output wire auto_bus_xing_in_d_bits_sink;
	output wire auto_bus_xing_in_d_bits_denied;
	output wire [31:0] auto_bus_xing_in_d_bits_data;
	output wire auto_bus_xing_in_d_bits_corrupt;
	input custom_boot;
	output wire clock;
	output wire reset;
	wire subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_clock;
	wire subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_reset;
	wire subsystem_cbus_clock_groups_auto_out_member_subsystem_cbus_0_clock;
	wire subsystem_cbus_clock_groups_auto_out_member_subsystem_cbus_0_reset;
	wire clockGroup_auto_in_member_subsystem_cbus_0_clock;
	wire clockGroup_auto_in_member_subsystem_cbus_0_reset;
	wire clockGroup_auto_out_clock;
	wire clockGroup_auto_out_reset;
	wire fixedClockNode_auto_in_clock;
	wire fixedClockNode_auto_in_reset;
	wire fixedClockNode_auto_out_5_clock;
	wire fixedClockNode_auto_out_5_reset;
	wire fixedClockNode_auto_out_4_clock;
	wire fixedClockNode_auto_out_4_reset;
	wire fixedClockNode_auto_out_3_clock;
	wire fixedClockNode_auto_out_3_reset;
	wire fixedClockNode_auto_out_1_clock;
	wire fixedClockNode_auto_out_1_reset;
	wire fixedClockNode_auto_out_0_clock;
	wire fixedClockNode_auto_out_0_reset;
	wire fixer_clock;
	wire fixer_reset;
	wire fixer_auto_in_a_ready;
	wire fixer_auto_in_a_valid;
	wire [2:0] fixer_auto_in_a_bits_opcode;
	wire [2:0] fixer_auto_in_a_bits_param;
	wire [3:0] fixer_auto_in_a_bits_size;
	wire [2:0] fixer_auto_in_a_bits_source;
	wire [31:0] fixer_auto_in_a_bits_address;
	wire [3:0] fixer_auto_in_a_bits_mask;
	wire [31:0] fixer_auto_in_a_bits_data;
	wire fixer_auto_in_a_bits_corrupt;
	wire fixer_auto_in_d_ready;
	wire fixer_auto_in_d_valid;
	wire [2:0] fixer_auto_in_d_bits_opcode;
	wire [1:0] fixer_auto_in_d_bits_param;
	wire [3:0] fixer_auto_in_d_bits_size;
	wire [2:0] fixer_auto_in_d_bits_source;
	wire fixer_auto_in_d_bits_sink;
	wire fixer_auto_in_d_bits_denied;
	wire [31:0] fixer_auto_in_d_bits_data;
	wire fixer_auto_in_d_bits_corrupt;
	wire fixer_auto_out_a_ready;
	wire fixer_auto_out_a_valid;
	wire [2:0] fixer_auto_out_a_bits_opcode;
	wire [2:0] fixer_auto_out_a_bits_param;
	wire [3:0] fixer_auto_out_a_bits_size;
	wire [2:0] fixer_auto_out_a_bits_source;
	wire [31:0] fixer_auto_out_a_bits_address;
	wire [3:0] fixer_auto_out_a_bits_mask;
	wire [31:0] fixer_auto_out_a_bits_data;
	wire fixer_auto_out_a_bits_corrupt;
	wire fixer_auto_out_d_ready;
	wire fixer_auto_out_d_valid;
	wire [2:0] fixer_auto_out_d_bits_opcode;
	wire [1:0] fixer_auto_out_d_bits_param;
	wire [3:0] fixer_auto_out_d_bits_size;
	wire [2:0] fixer_auto_out_d_bits_source;
	wire fixer_auto_out_d_bits_sink;
	wire fixer_auto_out_d_bits_denied;
	wire [31:0] fixer_auto_out_d_bits_data;
	wire fixer_auto_out_d_bits_corrupt;
	wire in_xbar_clock;
	wire in_xbar_reset;
	wire in_xbar_auto_in_1_a_ready;
	wire in_xbar_auto_in_1_a_valid;
	wire [31:0] in_xbar_auto_in_1_a_bits_address;
	wire [31:0] in_xbar_auto_in_1_a_bits_data;
	wire in_xbar_auto_in_1_d_valid;
	wire in_xbar_auto_in_0_a_ready;
	wire in_xbar_auto_in_0_a_valid;
	wire [2:0] in_xbar_auto_in_0_a_bits_opcode;
	wire [2:0] in_xbar_auto_in_0_a_bits_param;
	wire [3:0] in_xbar_auto_in_0_a_bits_size;
	wire [1:0] in_xbar_auto_in_0_a_bits_source;
	wire [31:0] in_xbar_auto_in_0_a_bits_address;
	wire [3:0] in_xbar_auto_in_0_a_bits_mask;
	wire [31:0] in_xbar_auto_in_0_a_bits_data;
	wire in_xbar_auto_in_0_a_bits_corrupt;
	wire in_xbar_auto_in_0_d_ready;
	wire in_xbar_auto_in_0_d_valid;
	wire [2:0] in_xbar_auto_in_0_d_bits_opcode;
	wire [1:0] in_xbar_auto_in_0_d_bits_param;
	wire [3:0] in_xbar_auto_in_0_d_bits_size;
	wire [1:0] in_xbar_auto_in_0_d_bits_source;
	wire in_xbar_auto_in_0_d_bits_sink;
	wire in_xbar_auto_in_0_d_bits_denied;
	wire [31:0] in_xbar_auto_in_0_d_bits_data;
	wire in_xbar_auto_in_0_d_bits_corrupt;
	wire in_xbar_auto_out_a_ready;
	wire in_xbar_auto_out_a_valid;
	wire [2:0] in_xbar_auto_out_a_bits_opcode;
	wire [2:0] in_xbar_auto_out_a_bits_param;
	wire [3:0] in_xbar_auto_out_a_bits_size;
	wire [2:0] in_xbar_auto_out_a_bits_source;
	wire [31:0] in_xbar_auto_out_a_bits_address;
	wire [3:0] in_xbar_auto_out_a_bits_mask;
	wire [31:0] in_xbar_auto_out_a_bits_data;
	wire in_xbar_auto_out_a_bits_corrupt;
	wire in_xbar_auto_out_d_ready;
	wire in_xbar_auto_out_d_valid;
	wire [2:0] in_xbar_auto_out_d_bits_opcode;
	wire [1:0] in_xbar_auto_out_d_bits_param;
	wire [3:0] in_xbar_auto_out_d_bits_size;
	wire [2:0] in_xbar_auto_out_d_bits_source;
	wire in_xbar_auto_out_d_bits_sink;
	wire in_xbar_auto_out_d_bits_denied;
	wire [31:0] in_xbar_auto_out_d_bits_data;
	wire in_xbar_auto_out_d_bits_corrupt;
	wire out_xbar_clock;
	wire out_xbar_reset;
	wire out_xbar_auto_in_a_ready;
	wire out_xbar_auto_in_a_valid;
	wire [2:0] out_xbar_auto_in_a_bits_opcode;
	wire [2:0] out_xbar_auto_in_a_bits_param;
	wire [3:0] out_xbar_auto_in_a_bits_size;
	wire [2:0] out_xbar_auto_in_a_bits_source;
	wire [31:0] out_xbar_auto_in_a_bits_address;
	wire [3:0] out_xbar_auto_in_a_bits_mask;
	wire [31:0] out_xbar_auto_in_a_bits_data;
	wire out_xbar_auto_in_a_bits_corrupt;
	wire out_xbar_auto_in_d_ready;
	wire out_xbar_auto_in_d_valid;
	wire [2:0] out_xbar_auto_in_d_bits_opcode;
	wire [1:0] out_xbar_auto_in_d_bits_param;
	wire [3:0] out_xbar_auto_in_d_bits_size;
	wire [2:0] out_xbar_auto_in_d_bits_source;
	wire out_xbar_auto_in_d_bits_sink;
	wire out_xbar_auto_in_d_bits_denied;
	wire [31:0] out_xbar_auto_in_d_bits_data;
	wire out_xbar_auto_in_d_bits_corrupt;
	wire out_xbar_auto_out_8_a_ready;
	wire out_xbar_auto_out_8_a_valid;
	wire [2:0] out_xbar_auto_out_8_a_bits_opcode;
	wire [2:0] out_xbar_auto_out_8_a_bits_param;
	wire [2:0] out_xbar_auto_out_8_a_bits_size;
	wire [2:0] out_xbar_auto_out_8_a_bits_source;
	wire [20:0] out_xbar_auto_out_8_a_bits_address;
	wire [3:0] out_xbar_auto_out_8_a_bits_mask;
	wire [31:0] out_xbar_auto_out_8_a_bits_data;
	wire out_xbar_auto_out_8_a_bits_corrupt;
	wire out_xbar_auto_out_8_d_ready;
	wire out_xbar_auto_out_8_d_valid;
	wire [2:0] out_xbar_auto_out_8_d_bits_opcode;
	wire [1:0] out_xbar_auto_out_8_d_bits_param;
	wire [2:0] out_xbar_auto_out_8_d_bits_size;
	wire [2:0] out_xbar_auto_out_8_d_bits_source;
	wire out_xbar_auto_out_8_d_bits_sink;
	wire out_xbar_auto_out_8_d_bits_denied;
	wire [31:0] out_xbar_auto_out_8_d_bits_data;
	wire out_xbar_auto_out_8_d_bits_corrupt;
	wire out_xbar_auto_out_7_a_ready;
	wire out_xbar_auto_out_7_a_valid;
	wire [2:0] out_xbar_auto_out_7_a_bits_opcode;
	wire [2:0] out_xbar_auto_out_7_a_bits_param;
	wire [2:0] out_xbar_auto_out_7_a_bits_size;
	wire [2:0] out_xbar_auto_out_7_a_bits_source;
	wire [20:0] out_xbar_auto_out_7_a_bits_address;
	wire [3:0] out_xbar_auto_out_7_a_bits_mask;
	wire [31:0] out_xbar_auto_out_7_a_bits_data;
	wire out_xbar_auto_out_7_a_bits_corrupt;
	wire out_xbar_auto_out_7_d_ready;
	wire out_xbar_auto_out_7_d_valid;
	wire [2:0] out_xbar_auto_out_7_d_bits_opcode;
	wire [1:0] out_xbar_auto_out_7_d_bits_param;
	wire [2:0] out_xbar_auto_out_7_d_bits_size;
	wire [2:0] out_xbar_auto_out_7_d_bits_source;
	wire out_xbar_auto_out_7_d_bits_sink;
	wire out_xbar_auto_out_7_d_bits_denied;
	wire [31:0] out_xbar_auto_out_7_d_bits_data;
	wire out_xbar_auto_out_7_d_bits_corrupt;
	wire out_xbar_auto_out_6_a_ready;
	wire out_xbar_auto_out_6_a_valid;
	wire [2:0] out_xbar_auto_out_6_a_bits_opcode;
	wire [2:0] out_xbar_auto_out_6_a_bits_param;
	wire [2:0] out_xbar_auto_out_6_a_bits_size;
	wire [2:0] out_xbar_auto_out_6_a_bits_source;
	wire [16:0] out_xbar_auto_out_6_a_bits_address;
	wire [3:0] out_xbar_auto_out_6_a_bits_mask;
	wire out_xbar_auto_out_6_a_bits_corrupt;
	wire out_xbar_auto_out_6_d_ready;
	wire out_xbar_auto_out_6_d_valid;
	wire [2:0] out_xbar_auto_out_6_d_bits_size;
	wire [2:0] out_xbar_auto_out_6_d_bits_source;
	wire [31:0] out_xbar_auto_out_6_d_bits_data;
	wire out_xbar_auto_out_5_a_ready;
	wire out_xbar_auto_out_5_a_valid;
	wire [2:0] out_xbar_auto_out_5_a_bits_opcode;
	wire [2:0] out_xbar_auto_out_5_a_bits_param;
	wire [2:0] out_xbar_auto_out_5_a_bits_size;
	wire [2:0] out_xbar_auto_out_5_a_bits_source;
	wire [31:0] out_xbar_auto_out_5_a_bits_address;
	wire [3:0] out_xbar_auto_out_5_a_bits_mask;
	wire [31:0] out_xbar_auto_out_5_a_bits_data;
	wire out_xbar_auto_out_5_d_ready;
	wire out_xbar_auto_out_5_d_valid;
	wire [2:0] out_xbar_auto_out_5_d_bits_opcode;
	wire [1:0] out_xbar_auto_out_5_d_bits_param;
	wire [2:0] out_xbar_auto_out_5_d_bits_size;
	wire [2:0] out_xbar_auto_out_5_d_bits_source;
	wire out_xbar_auto_out_5_d_bits_sink;
	wire out_xbar_auto_out_5_d_bits_denied;
	wire [31:0] out_xbar_auto_out_5_d_bits_data;
	wire out_xbar_auto_out_5_d_bits_corrupt;
	wire out_xbar_auto_out_4_a_ready;
	wire out_xbar_auto_out_4_a_valid;
	wire [2:0] out_xbar_auto_out_4_a_bits_opcode;
	wire [2:0] out_xbar_auto_out_4_a_bits_param;
	wire [2:0] out_xbar_auto_out_4_a_bits_size;
	wire [2:0] out_xbar_auto_out_4_a_bits_source;
	wire [11:0] out_xbar_auto_out_4_a_bits_address;
	wire [3:0] out_xbar_auto_out_4_a_bits_mask;
	wire [31:0] out_xbar_auto_out_4_a_bits_data;
	wire out_xbar_auto_out_4_a_bits_corrupt;
	wire out_xbar_auto_out_4_d_ready;
	wire out_xbar_auto_out_4_d_valid;
	wire [2:0] out_xbar_auto_out_4_d_bits_opcode;
	wire [2:0] out_xbar_auto_out_4_d_bits_size;
	wire [2:0] out_xbar_auto_out_4_d_bits_source;
	wire [31:0] out_xbar_auto_out_4_d_bits_data;
	wire out_xbar_auto_out_3_a_ready;
	wire out_xbar_auto_out_3_a_valid;
	wire [2:0] out_xbar_auto_out_3_a_bits_opcode;
	wire [2:0] out_xbar_auto_out_3_a_bits_param;
	wire [2:0] out_xbar_auto_out_3_a_bits_size;
	wire [2:0] out_xbar_auto_out_3_a_bits_source;
	wire [25:0] out_xbar_auto_out_3_a_bits_address;
	wire [3:0] out_xbar_auto_out_3_a_bits_mask;
	wire [31:0] out_xbar_auto_out_3_a_bits_data;
	wire out_xbar_auto_out_3_a_bits_corrupt;
	wire out_xbar_auto_out_3_d_ready;
	wire out_xbar_auto_out_3_d_valid;
	wire [2:0] out_xbar_auto_out_3_d_bits_opcode;
	wire [2:0] out_xbar_auto_out_3_d_bits_size;
	wire [2:0] out_xbar_auto_out_3_d_bits_source;
	wire [31:0] out_xbar_auto_out_3_d_bits_data;
	wire out_xbar_auto_out_2_a_ready;
	wire out_xbar_auto_out_2_a_valid;
	wire [2:0] out_xbar_auto_out_2_a_bits_opcode;
	wire [2:0] out_xbar_auto_out_2_a_bits_param;
	wire [2:0] out_xbar_auto_out_2_a_bits_size;
	wire [2:0] out_xbar_auto_out_2_a_bits_source;
	wire [27:0] out_xbar_auto_out_2_a_bits_address;
	wire [3:0] out_xbar_auto_out_2_a_bits_mask;
	wire [31:0] out_xbar_auto_out_2_a_bits_data;
	wire out_xbar_auto_out_2_a_bits_corrupt;
	wire out_xbar_auto_out_2_d_ready;
	wire out_xbar_auto_out_2_d_valid;
	wire [2:0] out_xbar_auto_out_2_d_bits_opcode;
	wire [2:0] out_xbar_auto_out_2_d_bits_size;
	wire [2:0] out_xbar_auto_out_2_d_bits_source;
	wire [31:0] out_xbar_auto_out_2_d_bits_data;
	wire out_xbar_auto_out_1_a_ready;
	wire out_xbar_auto_out_1_a_valid;
	wire [2:0] out_xbar_auto_out_1_a_bits_opcode;
	wire [2:0] out_xbar_auto_out_1_a_bits_param;
	wire [2:0] out_xbar_auto_out_1_a_bits_size;
	wire [2:0] out_xbar_auto_out_1_a_bits_source;
	wire [30:0] out_xbar_auto_out_1_a_bits_address;
	wire [3:0] out_xbar_auto_out_1_a_bits_mask;
	wire [31:0] out_xbar_auto_out_1_a_bits_data;
	wire out_xbar_auto_out_1_a_bits_corrupt;
	wire out_xbar_auto_out_1_d_ready;
	wire out_xbar_auto_out_1_d_valid;
	wire [2:0] out_xbar_auto_out_1_d_bits_opcode;
	wire [1:0] out_xbar_auto_out_1_d_bits_param;
	wire [2:0] out_xbar_auto_out_1_d_bits_size;
	wire [2:0] out_xbar_auto_out_1_d_bits_source;
	wire out_xbar_auto_out_1_d_bits_sink;
	wire out_xbar_auto_out_1_d_bits_denied;
	wire [31:0] out_xbar_auto_out_1_d_bits_data;
	wire out_xbar_auto_out_1_d_bits_corrupt;
	wire out_xbar_auto_out_0_a_ready;
	wire out_xbar_auto_out_0_a_valid;
	wire [2:0] out_xbar_auto_out_0_a_bits_opcode;
	wire [2:0] out_xbar_auto_out_0_a_bits_param;
	wire [3:0] out_xbar_auto_out_0_a_bits_size;
	wire [2:0] out_xbar_auto_out_0_a_bits_source;
	wire [13:0] out_xbar_auto_out_0_a_bits_address;
	wire [3:0] out_xbar_auto_out_0_a_bits_mask;
	wire out_xbar_auto_out_0_a_bits_corrupt;
	wire out_xbar_auto_out_0_d_ready;
	wire out_xbar_auto_out_0_d_valid;
	wire [2:0] out_xbar_auto_out_0_d_bits_opcode;
	wire [1:0] out_xbar_auto_out_0_d_bits_param;
	wire [3:0] out_xbar_auto_out_0_d_bits_size;
	wire [2:0] out_xbar_auto_out_0_d_bits_source;
	wire out_xbar_auto_out_0_d_bits_sink;
	wire out_xbar_auto_out_0_d_bits_denied;
	wire [31:0] out_xbar_auto_out_0_d_bits_data;
	wire out_xbar_auto_out_0_d_bits_corrupt;
	wire buffer_clock;
	wire buffer_reset;
	wire buffer_auto_in_a_ready;
	wire buffer_auto_in_a_valid;
	wire [2:0] buffer_auto_in_a_bits_opcode;
	wire [2:0] buffer_auto_in_a_bits_param;
	wire [3:0] buffer_auto_in_a_bits_size;
	wire [2:0] buffer_auto_in_a_bits_source;
	wire [31:0] buffer_auto_in_a_bits_address;
	wire [3:0] buffer_auto_in_a_bits_mask;
	wire [31:0] buffer_auto_in_a_bits_data;
	wire buffer_auto_in_a_bits_corrupt;
	wire buffer_auto_in_d_ready;
	wire buffer_auto_in_d_valid;
	wire [2:0] buffer_auto_in_d_bits_opcode;
	wire [1:0] buffer_auto_in_d_bits_param;
	wire [3:0] buffer_auto_in_d_bits_size;
	wire [2:0] buffer_auto_in_d_bits_source;
	wire buffer_auto_in_d_bits_sink;
	wire buffer_auto_in_d_bits_denied;
	wire [31:0] buffer_auto_in_d_bits_data;
	wire buffer_auto_in_d_bits_corrupt;
	wire buffer_auto_out_a_ready;
	wire buffer_auto_out_a_valid;
	wire [2:0] buffer_auto_out_a_bits_opcode;
	wire [2:0] buffer_auto_out_a_bits_param;
	wire [3:0] buffer_auto_out_a_bits_size;
	wire [2:0] buffer_auto_out_a_bits_source;
	wire [31:0] buffer_auto_out_a_bits_address;
	wire [3:0] buffer_auto_out_a_bits_mask;
	wire [31:0] buffer_auto_out_a_bits_data;
	wire buffer_auto_out_a_bits_corrupt;
	wire buffer_auto_out_d_ready;
	wire buffer_auto_out_d_valid;
	wire [2:0] buffer_auto_out_d_bits_opcode;
	wire [1:0] buffer_auto_out_d_bits_param;
	wire [3:0] buffer_auto_out_d_bits_size;
	wire [2:0] buffer_auto_out_d_bits_source;
	wire buffer_auto_out_d_bits_sink;
	wire buffer_auto_out_d_bits_denied;
	wire [31:0] buffer_auto_out_d_bits_data;
	wire buffer_auto_out_d_bits_corrupt;
	wire atomics_clock;
	wire atomics_reset;
	wire atomics_auto_in_a_ready;
	wire atomics_auto_in_a_valid;
	wire [2:0] atomics_auto_in_a_bits_opcode;
	wire [2:0] atomics_auto_in_a_bits_param;
	wire [3:0] atomics_auto_in_a_bits_size;
	wire [2:0] atomics_auto_in_a_bits_source;
	wire [31:0] atomics_auto_in_a_bits_address;
	wire [3:0] atomics_auto_in_a_bits_mask;
	wire [31:0] atomics_auto_in_a_bits_data;
	wire atomics_auto_in_a_bits_corrupt;
	wire atomics_auto_in_d_ready;
	wire atomics_auto_in_d_valid;
	wire [2:0] atomics_auto_in_d_bits_opcode;
	wire [1:0] atomics_auto_in_d_bits_param;
	wire [3:0] atomics_auto_in_d_bits_size;
	wire [2:0] atomics_auto_in_d_bits_source;
	wire atomics_auto_in_d_bits_sink;
	wire atomics_auto_in_d_bits_denied;
	wire [31:0] atomics_auto_in_d_bits_data;
	wire atomics_auto_in_d_bits_corrupt;
	wire atomics_auto_out_a_ready;
	wire atomics_auto_out_a_valid;
	wire [2:0] atomics_auto_out_a_bits_opcode;
	wire [2:0] atomics_auto_out_a_bits_param;
	wire [3:0] atomics_auto_out_a_bits_size;
	wire [2:0] atomics_auto_out_a_bits_source;
	wire [31:0] atomics_auto_out_a_bits_address;
	wire [3:0] atomics_auto_out_a_bits_mask;
	wire [31:0] atomics_auto_out_a_bits_data;
	wire atomics_auto_out_a_bits_corrupt;
	wire atomics_auto_out_d_ready;
	wire atomics_auto_out_d_valid;
	wire [2:0] atomics_auto_out_d_bits_opcode;
	wire [1:0] atomics_auto_out_d_bits_param;
	wire [3:0] atomics_auto_out_d_bits_size;
	wire [2:0] atomics_auto_out_d_bits_source;
	wire atomics_auto_out_d_bits_sink;
	wire atomics_auto_out_d_bits_denied;
	wire [31:0] atomics_auto_out_d_bits_data;
	wire atomics_auto_out_d_bits_corrupt;
	wire wrapped_error_device_clock;
	wire wrapped_error_device_reset;
	wire wrapped_error_device_auto_buffer_in_a_ready;
	wire wrapped_error_device_auto_buffer_in_a_valid;
	wire [2:0] wrapped_error_device_auto_buffer_in_a_bits_opcode;
	wire [2:0] wrapped_error_device_auto_buffer_in_a_bits_param;
	wire [3:0] wrapped_error_device_auto_buffer_in_a_bits_size;
	wire [2:0] wrapped_error_device_auto_buffer_in_a_bits_source;
	wire [13:0] wrapped_error_device_auto_buffer_in_a_bits_address;
	wire [3:0] wrapped_error_device_auto_buffer_in_a_bits_mask;
	wire wrapped_error_device_auto_buffer_in_a_bits_corrupt;
	wire wrapped_error_device_auto_buffer_in_d_ready;
	wire wrapped_error_device_auto_buffer_in_d_valid;
	wire [2:0] wrapped_error_device_auto_buffer_in_d_bits_opcode;
	wire [1:0] wrapped_error_device_auto_buffer_in_d_bits_param;
	wire [3:0] wrapped_error_device_auto_buffer_in_d_bits_size;
	wire [2:0] wrapped_error_device_auto_buffer_in_d_bits_source;
	wire wrapped_error_device_auto_buffer_in_d_bits_sink;
	wire wrapped_error_device_auto_buffer_in_d_bits_denied;
	wire [31:0] wrapped_error_device_auto_buffer_in_d_bits_data;
	wire wrapped_error_device_auto_buffer_in_d_bits_corrupt;
	wire buffer_1_auto_in_a_ready;
	wire buffer_1_auto_in_a_valid;
	wire [2:0] buffer_1_auto_in_a_bits_opcode;
	wire [2:0] buffer_1_auto_in_a_bits_param;
	wire [3:0] buffer_1_auto_in_a_bits_size;
	wire [1:0] buffer_1_auto_in_a_bits_source;
	wire [31:0] buffer_1_auto_in_a_bits_address;
	wire [3:0] buffer_1_auto_in_a_bits_mask;
	wire [31:0] buffer_1_auto_in_a_bits_data;
	wire buffer_1_auto_in_a_bits_corrupt;
	wire buffer_1_auto_in_d_ready;
	wire buffer_1_auto_in_d_valid;
	wire [2:0] buffer_1_auto_in_d_bits_opcode;
	wire [1:0] buffer_1_auto_in_d_bits_param;
	wire [3:0] buffer_1_auto_in_d_bits_size;
	wire [1:0] buffer_1_auto_in_d_bits_source;
	wire buffer_1_auto_in_d_bits_sink;
	wire buffer_1_auto_in_d_bits_denied;
	wire [31:0] buffer_1_auto_in_d_bits_data;
	wire buffer_1_auto_in_d_bits_corrupt;
	wire buffer_1_auto_out_a_ready;
	wire buffer_1_auto_out_a_valid;
	wire [2:0] buffer_1_auto_out_a_bits_opcode;
	wire [2:0] buffer_1_auto_out_a_bits_param;
	wire [3:0] buffer_1_auto_out_a_bits_size;
	wire [1:0] buffer_1_auto_out_a_bits_source;
	wire [31:0] buffer_1_auto_out_a_bits_address;
	wire [3:0] buffer_1_auto_out_a_bits_mask;
	wire [31:0] buffer_1_auto_out_a_bits_data;
	wire buffer_1_auto_out_a_bits_corrupt;
	wire buffer_1_auto_out_d_ready;
	wire buffer_1_auto_out_d_valid;
	wire [2:0] buffer_1_auto_out_d_bits_opcode;
	wire [1:0] buffer_1_auto_out_d_bits_param;
	wire [3:0] buffer_1_auto_out_d_bits_size;
	wire [1:0] buffer_1_auto_out_d_bits_source;
	wire buffer_1_auto_out_d_bits_sink;
	wire buffer_1_auto_out_d_bits_denied;
	wire [31:0] buffer_1_auto_out_d_bits_data;
	wire buffer_1_auto_out_d_bits_corrupt;
	wire coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_ready;
	wire coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_valid;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_opcode;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_param;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_size;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_source;
	wire [30:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_address;
	wire [3:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_mask;
	wire [31:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_data;
	wire coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_corrupt;
	wire coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_ready;
	wire coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_valid;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_opcode;
	wire [1:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_param;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_size;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_source;
	wire coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_sink;
	wire coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_denied;
	wire [31:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_data;
	wire coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_corrupt;
	wire coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_ready;
	wire coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_valid;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_opcode;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_param;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_size;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_source;
	wire [30:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_address;
	wire [3:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_mask;
	wire [31:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_data;
	wire coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_corrupt;
	wire coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_ready;
	wire coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_valid;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_opcode;
	wire [1:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_param;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_size;
	wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_source;
	wire coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_sink;
	wire coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_denied;
	wire [31:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_data;
	wire coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_corrupt;
	wire coupler_to_plic_clock;
	wire coupler_to_plic_reset;
	wire coupler_to_plic_auto_fragmenter_out_a_ready;
	wire coupler_to_plic_auto_fragmenter_out_a_valid;
	wire [2:0] coupler_to_plic_auto_fragmenter_out_a_bits_opcode;
	wire [2:0] coupler_to_plic_auto_fragmenter_out_a_bits_param;
	wire [1:0] coupler_to_plic_auto_fragmenter_out_a_bits_size;
	wire [7:0] coupler_to_plic_auto_fragmenter_out_a_bits_source;
	wire [27:0] coupler_to_plic_auto_fragmenter_out_a_bits_address;
	wire [3:0] coupler_to_plic_auto_fragmenter_out_a_bits_mask;
	wire [31:0] coupler_to_plic_auto_fragmenter_out_a_bits_data;
	wire coupler_to_plic_auto_fragmenter_out_a_bits_corrupt;
	wire coupler_to_plic_auto_fragmenter_out_d_ready;
	wire coupler_to_plic_auto_fragmenter_out_d_valid;
	wire [2:0] coupler_to_plic_auto_fragmenter_out_d_bits_opcode;
	wire [1:0] coupler_to_plic_auto_fragmenter_out_d_bits_size;
	wire [7:0] coupler_to_plic_auto_fragmenter_out_d_bits_source;
	wire [31:0] coupler_to_plic_auto_fragmenter_out_d_bits_data;
	wire coupler_to_plic_auto_tl_in_a_ready;
	wire coupler_to_plic_auto_tl_in_a_valid;
	wire [2:0] coupler_to_plic_auto_tl_in_a_bits_opcode;
	wire [2:0] coupler_to_plic_auto_tl_in_a_bits_param;
	wire [2:0] coupler_to_plic_auto_tl_in_a_bits_size;
	wire [2:0] coupler_to_plic_auto_tl_in_a_bits_source;
	wire [27:0] coupler_to_plic_auto_tl_in_a_bits_address;
	wire [3:0] coupler_to_plic_auto_tl_in_a_bits_mask;
	wire [31:0] coupler_to_plic_auto_tl_in_a_bits_data;
	wire coupler_to_plic_auto_tl_in_a_bits_corrupt;
	wire coupler_to_plic_auto_tl_in_d_ready;
	wire coupler_to_plic_auto_tl_in_d_valid;
	wire [2:0] coupler_to_plic_auto_tl_in_d_bits_opcode;
	wire [2:0] coupler_to_plic_auto_tl_in_d_bits_size;
	wire [2:0] coupler_to_plic_auto_tl_in_d_bits_source;
	wire [31:0] coupler_to_plic_auto_tl_in_d_bits_data;
	wire coupler_to_clint_clock;
	wire coupler_to_clint_reset;
	wire coupler_to_clint_auto_fragmenter_out_a_ready;
	wire coupler_to_clint_auto_fragmenter_out_a_valid;
	wire [2:0] coupler_to_clint_auto_fragmenter_out_a_bits_opcode;
	wire [2:0] coupler_to_clint_auto_fragmenter_out_a_bits_param;
	wire [1:0] coupler_to_clint_auto_fragmenter_out_a_bits_size;
	wire [7:0] coupler_to_clint_auto_fragmenter_out_a_bits_source;
	wire [25:0] coupler_to_clint_auto_fragmenter_out_a_bits_address;
	wire [3:0] coupler_to_clint_auto_fragmenter_out_a_bits_mask;
	wire [31:0] coupler_to_clint_auto_fragmenter_out_a_bits_data;
	wire coupler_to_clint_auto_fragmenter_out_a_bits_corrupt;
	wire coupler_to_clint_auto_fragmenter_out_d_ready;
	wire coupler_to_clint_auto_fragmenter_out_d_valid;
	wire [2:0] coupler_to_clint_auto_fragmenter_out_d_bits_opcode;
	wire [1:0] coupler_to_clint_auto_fragmenter_out_d_bits_size;
	wire [7:0] coupler_to_clint_auto_fragmenter_out_d_bits_source;
	wire [31:0] coupler_to_clint_auto_fragmenter_out_d_bits_data;
	wire coupler_to_clint_auto_tl_in_a_ready;
	wire coupler_to_clint_auto_tl_in_a_valid;
	wire [2:0] coupler_to_clint_auto_tl_in_a_bits_opcode;
	wire [2:0] coupler_to_clint_auto_tl_in_a_bits_param;
	wire [2:0] coupler_to_clint_auto_tl_in_a_bits_size;
	wire [2:0] coupler_to_clint_auto_tl_in_a_bits_source;
	wire [25:0] coupler_to_clint_auto_tl_in_a_bits_address;
	wire [3:0] coupler_to_clint_auto_tl_in_a_bits_mask;
	wire [31:0] coupler_to_clint_auto_tl_in_a_bits_data;
	wire coupler_to_clint_auto_tl_in_a_bits_corrupt;
	wire coupler_to_clint_auto_tl_in_d_ready;
	wire coupler_to_clint_auto_tl_in_d_valid;
	wire [2:0] coupler_to_clint_auto_tl_in_d_bits_opcode;
	wire [2:0] coupler_to_clint_auto_tl_in_d_bits_size;
	wire [2:0] coupler_to_clint_auto_tl_in_d_bits_source;
	wire [31:0] coupler_to_clint_auto_tl_in_d_bits_data;
	wire coupler_to_debug_clock;
	wire coupler_to_debug_reset;
	wire coupler_to_debug_auto_fragmenter_out_a_ready;
	wire coupler_to_debug_auto_fragmenter_out_a_valid;
	wire [2:0] coupler_to_debug_auto_fragmenter_out_a_bits_opcode;
	wire [2:0] coupler_to_debug_auto_fragmenter_out_a_bits_param;
	wire [1:0] coupler_to_debug_auto_fragmenter_out_a_bits_size;
	wire [7:0] coupler_to_debug_auto_fragmenter_out_a_bits_source;
	wire [11:0] coupler_to_debug_auto_fragmenter_out_a_bits_address;
	wire [3:0] coupler_to_debug_auto_fragmenter_out_a_bits_mask;
	wire [31:0] coupler_to_debug_auto_fragmenter_out_a_bits_data;
	wire coupler_to_debug_auto_fragmenter_out_a_bits_corrupt;
	wire coupler_to_debug_auto_fragmenter_out_d_ready;
	wire coupler_to_debug_auto_fragmenter_out_d_valid;
	wire [2:0] coupler_to_debug_auto_fragmenter_out_d_bits_opcode;
	wire [1:0] coupler_to_debug_auto_fragmenter_out_d_bits_size;
	wire [7:0] coupler_to_debug_auto_fragmenter_out_d_bits_source;
	wire [31:0] coupler_to_debug_auto_fragmenter_out_d_bits_data;
	wire coupler_to_debug_auto_tl_in_a_ready;
	wire coupler_to_debug_auto_tl_in_a_valid;
	wire [2:0] coupler_to_debug_auto_tl_in_a_bits_opcode;
	wire [2:0] coupler_to_debug_auto_tl_in_a_bits_param;
	wire [2:0] coupler_to_debug_auto_tl_in_a_bits_size;
	wire [2:0] coupler_to_debug_auto_tl_in_a_bits_source;
	wire [11:0] coupler_to_debug_auto_tl_in_a_bits_address;
	wire [3:0] coupler_to_debug_auto_tl_in_a_bits_mask;
	wire [31:0] coupler_to_debug_auto_tl_in_a_bits_data;
	wire coupler_to_debug_auto_tl_in_a_bits_corrupt;
	wire coupler_to_debug_auto_tl_in_d_ready;
	wire coupler_to_debug_auto_tl_in_d_valid;
	wire [2:0] coupler_to_debug_auto_tl_in_d_bits_opcode;
	wire [2:0] coupler_to_debug_auto_tl_in_d_bits_size;
	wire [2:0] coupler_to_debug_auto_tl_in_d_bits_source;
	wire [31:0] coupler_to_debug_auto_tl_in_d_bits_data;
	wire coupler_to_tile_auto_tl_slave_clock_xing_out_a_ready;
	wire coupler_to_tile_auto_tl_slave_clock_xing_out_a_valid;
	wire [2:0] coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_opcode;
	wire [2:0] coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_param;
	wire [2:0] coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_size;
	wire [2:0] coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_source;
	wire [31:0] coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_address;
	wire [3:0] coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_mask;
	wire [31:0] coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_data;
	wire coupler_to_tile_auto_tl_slave_clock_xing_out_d_ready;
	wire coupler_to_tile_auto_tl_slave_clock_xing_out_d_valid;
	wire [2:0] coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_opcode;
	wire [1:0] coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_param;
	wire [2:0] coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_size;
	wire [2:0] coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_source;
	wire coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_sink;
	wire coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_denied;
	wire [31:0] coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_data;
	wire coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_corrupt;
	wire coupler_to_tile_auto_tl_in_a_ready;
	wire coupler_to_tile_auto_tl_in_a_valid;
	wire [2:0] coupler_to_tile_auto_tl_in_a_bits_opcode;
	wire [2:0] coupler_to_tile_auto_tl_in_a_bits_param;
	wire [2:0] coupler_to_tile_auto_tl_in_a_bits_size;
	wire [2:0] coupler_to_tile_auto_tl_in_a_bits_source;
	wire [31:0] coupler_to_tile_auto_tl_in_a_bits_address;
	wire [3:0] coupler_to_tile_auto_tl_in_a_bits_mask;
	wire [31:0] coupler_to_tile_auto_tl_in_a_bits_data;
	wire coupler_to_tile_auto_tl_in_d_ready;
	wire coupler_to_tile_auto_tl_in_d_valid;
	wire [2:0] coupler_to_tile_auto_tl_in_d_bits_opcode;
	wire [1:0] coupler_to_tile_auto_tl_in_d_bits_param;
	wire [2:0] coupler_to_tile_auto_tl_in_d_bits_size;
	wire [2:0] coupler_to_tile_auto_tl_in_d_bits_source;
	wire coupler_to_tile_auto_tl_in_d_bits_sink;
	wire coupler_to_tile_auto_tl_in_d_bits_denied;
	wire [31:0] coupler_to_tile_auto_tl_in_d_bits_data;
	wire coupler_to_tile_auto_tl_in_d_bits_corrupt;
	wire coupler_to_bootrom_clock;
	wire coupler_to_bootrom_reset;
	wire coupler_to_bootrom_auto_fragmenter_out_a_ready;
	wire coupler_to_bootrom_auto_fragmenter_out_a_valid;
	wire [2:0] coupler_to_bootrom_auto_fragmenter_out_a_bits_opcode;
	wire [2:0] coupler_to_bootrom_auto_fragmenter_out_a_bits_param;
	wire [1:0] coupler_to_bootrom_auto_fragmenter_out_a_bits_size;
	wire [7:0] coupler_to_bootrom_auto_fragmenter_out_a_bits_source;
	wire [16:0] coupler_to_bootrom_auto_fragmenter_out_a_bits_address;
	wire [3:0] coupler_to_bootrom_auto_fragmenter_out_a_bits_mask;
	wire coupler_to_bootrom_auto_fragmenter_out_a_bits_corrupt;
	wire coupler_to_bootrom_auto_fragmenter_out_d_ready;
	wire coupler_to_bootrom_auto_fragmenter_out_d_valid;
	wire [1:0] coupler_to_bootrom_auto_fragmenter_out_d_bits_size;
	wire [7:0] coupler_to_bootrom_auto_fragmenter_out_d_bits_source;
	wire [31:0] coupler_to_bootrom_auto_fragmenter_out_d_bits_data;
	wire coupler_to_bootrom_auto_tl_in_a_ready;
	wire coupler_to_bootrom_auto_tl_in_a_valid;
	wire [2:0] coupler_to_bootrom_auto_tl_in_a_bits_opcode;
	wire [2:0] coupler_to_bootrom_auto_tl_in_a_bits_param;
	wire [2:0] coupler_to_bootrom_auto_tl_in_a_bits_size;
	wire [2:0] coupler_to_bootrom_auto_tl_in_a_bits_source;
	wire [16:0] coupler_to_bootrom_auto_tl_in_a_bits_address;
	wire [3:0] coupler_to_bootrom_auto_tl_in_a_bits_mask;
	wire coupler_to_bootrom_auto_tl_in_a_bits_corrupt;
	wire coupler_to_bootrom_auto_tl_in_d_ready;
	wire coupler_to_bootrom_auto_tl_in_d_valid;
	wire [2:0] coupler_to_bootrom_auto_tl_in_d_bits_size;
	wire [2:0] coupler_to_bootrom_auto_tl_in_d_bits_source;
	wire [31:0] coupler_to_bootrom_auto_tl_in_d_bits_data;
	wire coupler_from_port_named_custom_boot_pin_auto_tl_in_a_ready;
	wire coupler_from_port_named_custom_boot_pin_auto_tl_in_a_valid;
	wire [31:0] coupler_from_port_named_custom_boot_pin_auto_tl_in_a_bits_address;
	wire [31:0] coupler_from_port_named_custom_boot_pin_auto_tl_in_a_bits_data;
	wire coupler_from_port_named_custom_boot_pin_auto_tl_in_d_valid;
	wire coupler_from_port_named_custom_boot_pin_auto_tl_out_a_ready;
	wire coupler_from_port_named_custom_boot_pin_auto_tl_out_a_valid;
	wire [31:0] coupler_from_port_named_custom_boot_pin_auto_tl_out_a_bits_address;
	wire [31:0] coupler_from_port_named_custom_boot_pin_auto_tl_out_a_bits_data;
	wire coupler_from_port_named_custom_boot_pin_auto_tl_out_d_valid;
	wire coupler_to_slave_named_clockgater_clock;
	wire coupler_to_slave_named_clockgater_reset;
	wire coupler_to_slave_named_clockgater_auto_buffer_in_a_ready;
	wire coupler_to_slave_named_clockgater_auto_buffer_in_a_valid;
	wire [2:0] coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_opcode;
	wire [2:0] coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_param;
	wire [2:0] coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_size;
	wire [2:0] coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_source;
	wire [20:0] coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_address;
	wire [3:0] coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_mask;
	wire [31:0] coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_data;
	wire coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_corrupt;
	wire coupler_to_slave_named_clockgater_auto_buffer_in_d_ready;
	wire coupler_to_slave_named_clockgater_auto_buffer_in_d_valid;
	wire [2:0] coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_opcode;
	wire [1:0] coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_param;
	wire [2:0] coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_size;
	wire [2:0] coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_source;
	wire coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_sink;
	wire coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_denied;
	wire [31:0] coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_data;
	wire coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_corrupt;
	wire coupler_to_slave_named_clockgater_auto_buffer_out_a_ready;
	wire coupler_to_slave_named_clockgater_auto_buffer_out_a_valid;
	wire [2:0] coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_opcode;
	wire [2:0] coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_param;
	wire [1:0] coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_size;
	wire [7:0] coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_source;
	wire [20:0] coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_address;
	wire [3:0] coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_mask;
	wire [31:0] coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_data;
	wire coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_corrupt;
	wire coupler_to_slave_named_clockgater_auto_buffer_out_d_ready;
	wire coupler_to_slave_named_clockgater_auto_buffer_out_d_valid;
	wire [2:0] coupler_to_slave_named_clockgater_auto_buffer_out_d_bits_opcode;
	wire [1:0] coupler_to_slave_named_clockgater_auto_buffer_out_d_bits_size;
	wire [7:0] coupler_to_slave_named_clockgater_auto_buffer_out_d_bits_source;
	wire [31:0] coupler_to_slave_named_clockgater_auto_buffer_out_d_bits_data;
	wire coupler_to_slave_named_tileresetsetter_clock;
	wire coupler_to_slave_named_tileresetsetter_reset;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_ready;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_valid;
	wire [2:0] coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_opcode;
	wire [2:0] coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_param;
	wire [2:0] coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_size;
	wire [2:0] coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_source;
	wire [20:0] coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_address;
	wire [3:0] coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_mask;
	wire [31:0] coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_data;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_corrupt;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_ready;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_valid;
	wire [2:0] coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_opcode;
	wire [1:0] coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_param;
	wire [2:0] coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_size;
	wire [2:0] coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_source;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_sink;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_denied;
	wire [31:0] coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_data;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_corrupt;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_ready;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_valid;
	wire [2:0] coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_opcode;
	wire [2:0] coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_param;
	wire [1:0] coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_size;
	wire [7:0] coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_source;
	wire [20:0] coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_address;
	wire [3:0] coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_mask;
	wire [31:0] coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_data;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_corrupt;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_ready;
	wire coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_valid;
	wire [2:0] coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_bits_opcode;
	wire [1:0] coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_bits_size;
	wire [7:0] coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_bits_source;
	wire [31:0] coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_bits_data;
	wire bundleIn_0_clock = fixedClockNode_auto_out_0_clock;
	reg [2:0] state;
	wire bundleOut_0_1_a_ready = coupler_from_port_named_custom_boot_pin_auto_tl_in_a_ready;
	wire _GEN_19 = (3'h2 == state ? 1'h0 : 3'h3 == state);
	wire _GEN_28 = (3'h1 == state) | _GEN_19;
	wire bundleOut_0_1_a_valid = (3'h0 == state ? 1'h0 : _GEN_28);
	wire _T_2 = bundleOut_0_1_a_ready & bundleOut_0_1_a_valid;
	wire bundleOut_0_1_d_valid = coupler_from_port_named_custom_boot_pin_auto_tl_in_d_valid;
	wire [2:0] _GEN_2 = (bundleOut_0_1_d_valid ? 3'h3 : state);
	wire [2:0] _GEN_3 = (_T_2 ? 3'h4 : state);
	wire [2:0] _GEN_4 = (bundleOut_0_1_d_valid ? 3'h5 : state);
	wire [2:0] _GEN_5 = (~custom_boot ? 3'h0 : state);
	wire [2:0] _GEN_6 = (3'h5 == state ? _GEN_5 : state);
	wire [2:0] _GEN_7 = (3'h4 == state ? _GEN_4 : _GEN_6);
	wire [2:0] _GEN_17 = (3'h3 == state ? _GEN_3 : _GEN_7);
	wire bundleIn_0_reset = fixedClockNode_auto_out_0_reset;
	ClockGroupAggregator_3 subsystem_cbus_clock_groups(
		.auto_in_member_subsystem_cbus_0_clock(subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_clock),
		.auto_in_member_subsystem_cbus_0_reset(subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_reset),
		.auto_out_member_subsystem_cbus_0_clock(subsystem_cbus_clock_groups_auto_out_member_subsystem_cbus_0_clock),
		.auto_out_member_subsystem_cbus_0_reset(subsystem_cbus_clock_groups_auto_out_member_subsystem_cbus_0_reset)
	);
	ClockGroup_3 clockGroup(
		.auto_in_member_subsystem_cbus_0_clock(clockGroup_auto_in_member_subsystem_cbus_0_clock),
		.auto_in_member_subsystem_cbus_0_reset(clockGroup_auto_in_member_subsystem_cbus_0_reset),
		.auto_out_clock(clockGroup_auto_out_clock),
		.auto_out_reset(clockGroup_auto_out_reset)
	);
	FixedClockBroadcast_3 fixedClockNode(
		.auto_in_clock(fixedClockNode_auto_in_clock),
		.auto_in_reset(fixedClockNode_auto_in_reset),
		.auto_out_5_clock(fixedClockNode_auto_out_5_clock),
		.auto_out_5_reset(fixedClockNode_auto_out_5_reset),
		.auto_out_4_clock(fixedClockNode_auto_out_4_clock),
		.auto_out_4_reset(fixedClockNode_auto_out_4_reset),
		.auto_out_3_clock(fixedClockNode_auto_out_3_clock),
		.auto_out_3_reset(fixedClockNode_auto_out_3_reset),
		.auto_out_1_clock(fixedClockNode_auto_out_1_clock),
		.auto_out_1_reset(fixedClockNode_auto_out_1_reset),
		.auto_out_0_clock(fixedClockNode_auto_out_0_clock),
		.auto_out_0_reset(fixedClockNode_auto_out_0_reset)
	);
	TLFIFOFixer_2 fixer(
		.clock(fixer_clock),
		.reset(fixer_reset),
		.auto_in_a_ready(fixer_auto_in_a_ready),
		.auto_in_a_valid(fixer_auto_in_a_valid),
		.auto_in_a_bits_opcode(fixer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(fixer_auto_in_a_bits_param),
		.auto_in_a_bits_size(fixer_auto_in_a_bits_size),
		.auto_in_a_bits_source(fixer_auto_in_a_bits_source),
		.auto_in_a_bits_address(fixer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(fixer_auto_in_a_bits_mask),
		.auto_in_a_bits_data(fixer_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(fixer_auto_in_a_bits_corrupt),
		.auto_in_d_ready(fixer_auto_in_d_ready),
		.auto_in_d_valid(fixer_auto_in_d_valid),
		.auto_in_d_bits_opcode(fixer_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(fixer_auto_in_d_bits_param),
		.auto_in_d_bits_size(fixer_auto_in_d_bits_size),
		.auto_in_d_bits_source(fixer_auto_in_d_bits_source),
		.auto_in_d_bits_sink(fixer_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(fixer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(fixer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(fixer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(fixer_auto_out_a_ready),
		.auto_out_a_valid(fixer_auto_out_a_valid),
		.auto_out_a_bits_opcode(fixer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(fixer_auto_out_a_bits_param),
		.auto_out_a_bits_size(fixer_auto_out_a_bits_size),
		.auto_out_a_bits_source(fixer_auto_out_a_bits_source),
		.auto_out_a_bits_address(fixer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(fixer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(fixer_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(fixer_auto_out_a_bits_corrupt),
		.auto_out_d_ready(fixer_auto_out_d_ready),
		.auto_out_d_valid(fixer_auto_out_d_valid),
		.auto_out_d_bits_opcode(fixer_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(fixer_auto_out_d_bits_param),
		.auto_out_d_bits_size(fixer_auto_out_d_bits_size),
		.auto_out_d_bits_source(fixer_auto_out_d_bits_source),
		.auto_out_d_bits_sink(fixer_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(fixer_auto_out_d_bits_denied),
		.auto_out_d_bits_data(fixer_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(fixer_auto_out_d_bits_corrupt)
	);
	TLXbar_4 in_xbar(
		.clock(in_xbar_clock),
		.reset(in_xbar_reset),
		.auto_in_1_a_ready(in_xbar_auto_in_1_a_ready),
		.auto_in_1_a_valid(in_xbar_auto_in_1_a_valid),
		.auto_in_1_a_bits_address(in_xbar_auto_in_1_a_bits_address),
		.auto_in_1_a_bits_data(in_xbar_auto_in_1_a_bits_data),
		.auto_in_1_d_valid(in_xbar_auto_in_1_d_valid),
		.auto_in_0_a_ready(in_xbar_auto_in_0_a_ready),
		.auto_in_0_a_valid(in_xbar_auto_in_0_a_valid),
		.auto_in_0_a_bits_opcode(in_xbar_auto_in_0_a_bits_opcode),
		.auto_in_0_a_bits_param(in_xbar_auto_in_0_a_bits_param),
		.auto_in_0_a_bits_size(in_xbar_auto_in_0_a_bits_size),
		.auto_in_0_a_bits_source(in_xbar_auto_in_0_a_bits_source),
		.auto_in_0_a_bits_address(in_xbar_auto_in_0_a_bits_address),
		.auto_in_0_a_bits_mask(in_xbar_auto_in_0_a_bits_mask),
		.auto_in_0_a_bits_data(in_xbar_auto_in_0_a_bits_data),
		.auto_in_0_a_bits_corrupt(in_xbar_auto_in_0_a_bits_corrupt),
		.auto_in_0_d_ready(in_xbar_auto_in_0_d_ready),
		.auto_in_0_d_valid(in_xbar_auto_in_0_d_valid),
		.auto_in_0_d_bits_opcode(in_xbar_auto_in_0_d_bits_opcode),
		.auto_in_0_d_bits_param(in_xbar_auto_in_0_d_bits_param),
		.auto_in_0_d_bits_size(in_xbar_auto_in_0_d_bits_size),
		.auto_in_0_d_bits_source(in_xbar_auto_in_0_d_bits_source),
		.auto_in_0_d_bits_sink(in_xbar_auto_in_0_d_bits_sink),
		.auto_in_0_d_bits_denied(in_xbar_auto_in_0_d_bits_denied),
		.auto_in_0_d_bits_data(in_xbar_auto_in_0_d_bits_data),
		.auto_in_0_d_bits_corrupt(in_xbar_auto_in_0_d_bits_corrupt),
		.auto_out_a_ready(in_xbar_auto_out_a_ready),
		.auto_out_a_valid(in_xbar_auto_out_a_valid),
		.auto_out_a_bits_opcode(in_xbar_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(in_xbar_auto_out_a_bits_param),
		.auto_out_a_bits_size(in_xbar_auto_out_a_bits_size),
		.auto_out_a_bits_source(in_xbar_auto_out_a_bits_source),
		.auto_out_a_bits_address(in_xbar_auto_out_a_bits_address),
		.auto_out_a_bits_mask(in_xbar_auto_out_a_bits_mask),
		.auto_out_a_bits_data(in_xbar_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(in_xbar_auto_out_a_bits_corrupt),
		.auto_out_d_ready(in_xbar_auto_out_d_ready),
		.auto_out_d_valid(in_xbar_auto_out_d_valid),
		.auto_out_d_bits_opcode(in_xbar_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(in_xbar_auto_out_d_bits_param),
		.auto_out_d_bits_size(in_xbar_auto_out_d_bits_size),
		.auto_out_d_bits_source(in_xbar_auto_out_d_bits_source),
		.auto_out_d_bits_sink(in_xbar_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(in_xbar_auto_out_d_bits_denied),
		.auto_out_d_bits_data(in_xbar_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(in_xbar_auto_out_d_bits_corrupt)
	);
	TLXbar_5 out_xbar(
		.clock(out_xbar_clock),
		.reset(out_xbar_reset),
		.auto_in_a_ready(out_xbar_auto_in_a_ready),
		.auto_in_a_valid(out_xbar_auto_in_a_valid),
		.auto_in_a_bits_opcode(out_xbar_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(out_xbar_auto_in_a_bits_param),
		.auto_in_a_bits_size(out_xbar_auto_in_a_bits_size),
		.auto_in_a_bits_source(out_xbar_auto_in_a_bits_source),
		.auto_in_a_bits_address(out_xbar_auto_in_a_bits_address),
		.auto_in_a_bits_mask(out_xbar_auto_in_a_bits_mask),
		.auto_in_a_bits_data(out_xbar_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(out_xbar_auto_in_a_bits_corrupt),
		.auto_in_d_ready(out_xbar_auto_in_d_ready),
		.auto_in_d_valid(out_xbar_auto_in_d_valid),
		.auto_in_d_bits_opcode(out_xbar_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(out_xbar_auto_in_d_bits_param),
		.auto_in_d_bits_size(out_xbar_auto_in_d_bits_size),
		.auto_in_d_bits_source(out_xbar_auto_in_d_bits_source),
		.auto_in_d_bits_sink(out_xbar_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(out_xbar_auto_in_d_bits_denied),
		.auto_in_d_bits_data(out_xbar_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(out_xbar_auto_in_d_bits_corrupt),
		.auto_out_8_a_ready(out_xbar_auto_out_8_a_ready),
		.auto_out_8_a_valid(out_xbar_auto_out_8_a_valid),
		.auto_out_8_a_bits_opcode(out_xbar_auto_out_8_a_bits_opcode),
		.auto_out_8_a_bits_param(out_xbar_auto_out_8_a_bits_param),
		.auto_out_8_a_bits_size(out_xbar_auto_out_8_a_bits_size),
		.auto_out_8_a_bits_source(out_xbar_auto_out_8_a_bits_source),
		.auto_out_8_a_bits_address(out_xbar_auto_out_8_a_bits_address),
		.auto_out_8_a_bits_mask(out_xbar_auto_out_8_a_bits_mask),
		.auto_out_8_a_bits_data(out_xbar_auto_out_8_a_bits_data),
		.auto_out_8_a_bits_corrupt(out_xbar_auto_out_8_a_bits_corrupt),
		.auto_out_8_d_ready(out_xbar_auto_out_8_d_ready),
		.auto_out_8_d_valid(out_xbar_auto_out_8_d_valid),
		.auto_out_8_d_bits_opcode(out_xbar_auto_out_8_d_bits_opcode),
		.auto_out_8_d_bits_param(out_xbar_auto_out_8_d_bits_param),
		.auto_out_8_d_bits_size(out_xbar_auto_out_8_d_bits_size),
		.auto_out_8_d_bits_source(out_xbar_auto_out_8_d_bits_source),
		.auto_out_8_d_bits_sink(out_xbar_auto_out_8_d_bits_sink),
		.auto_out_8_d_bits_denied(out_xbar_auto_out_8_d_bits_denied),
		.auto_out_8_d_bits_data(out_xbar_auto_out_8_d_bits_data),
		.auto_out_8_d_bits_corrupt(out_xbar_auto_out_8_d_bits_corrupt),
		.auto_out_7_a_ready(out_xbar_auto_out_7_a_ready),
		.auto_out_7_a_valid(out_xbar_auto_out_7_a_valid),
		.auto_out_7_a_bits_opcode(out_xbar_auto_out_7_a_bits_opcode),
		.auto_out_7_a_bits_param(out_xbar_auto_out_7_a_bits_param),
		.auto_out_7_a_bits_size(out_xbar_auto_out_7_a_bits_size),
		.auto_out_7_a_bits_source(out_xbar_auto_out_7_a_bits_source),
		.auto_out_7_a_bits_address(out_xbar_auto_out_7_a_bits_address),
		.auto_out_7_a_bits_mask(out_xbar_auto_out_7_a_bits_mask),
		.auto_out_7_a_bits_data(out_xbar_auto_out_7_a_bits_data),
		.auto_out_7_a_bits_corrupt(out_xbar_auto_out_7_a_bits_corrupt),
		.auto_out_7_d_ready(out_xbar_auto_out_7_d_ready),
		.auto_out_7_d_valid(out_xbar_auto_out_7_d_valid),
		.auto_out_7_d_bits_opcode(out_xbar_auto_out_7_d_bits_opcode),
		.auto_out_7_d_bits_param(out_xbar_auto_out_7_d_bits_param),
		.auto_out_7_d_bits_size(out_xbar_auto_out_7_d_bits_size),
		.auto_out_7_d_bits_source(out_xbar_auto_out_7_d_bits_source),
		.auto_out_7_d_bits_sink(out_xbar_auto_out_7_d_bits_sink),
		.auto_out_7_d_bits_denied(out_xbar_auto_out_7_d_bits_denied),
		.auto_out_7_d_bits_data(out_xbar_auto_out_7_d_bits_data),
		.auto_out_7_d_bits_corrupt(out_xbar_auto_out_7_d_bits_corrupt),
		.auto_out_6_a_ready(out_xbar_auto_out_6_a_ready),
		.auto_out_6_a_valid(out_xbar_auto_out_6_a_valid),
		.auto_out_6_a_bits_opcode(out_xbar_auto_out_6_a_bits_opcode),
		.auto_out_6_a_bits_param(out_xbar_auto_out_6_a_bits_param),
		.auto_out_6_a_bits_size(out_xbar_auto_out_6_a_bits_size),
		.auto_out_6_a_bits_source(out_xbar_auto_out_6_a_bits_source),
		.auto_out_6_a_bits_address(out_xbar_auto_out_6_a_bits_address),
		.auto_out_6_a_bits_mask(out_xbar_auto_out_6_a_bits_mask),
		.auto_out_6_a_bits_corrupt(out_xbar_auto_out_6_a_bits_corrupt),
		.auto_out_6_d_ready(out_xbar_auto_out_6_d_ready),
		.auto_out_6_d_valid(out_xbar_auto_out_6_d_valid),
		.auto_out_6_d_bits_size(out_xbar_auto_out_6_d_bits_size),
		.auto_out_6_d_bits_source(out_xbar_auto_out_6_d_bits_source),
		.auto_out_6_d_bits_data(out_xbar_auto_out_6_d_bits_data),
		.auto_out_5_a_ready(out_xbar_auto_out_5_a_ready),
		.auto_out_5_a_valid(out_xbar_auto_out_5_a_valid),
		.auto_out_5_a_bits_opcode(out_xbar_auto_out_5_a_bits_opcode),
		.auto_out_5_a_bits_param(out_xbar_auto_out_5_a_bits_param),
		.auto_out_5_a_bits_size(out_xbar_auto_out_5_a_bits_size),
		.auto_out_5_a_bits_source(out_xbar_auto_out_5_a_bits_source),
		.auto_out_5_a_bits_address(out_xbar_auto_out_5_a_bits_address),
		.auto_out_5_a_bits_mask(out_xbar_auto_out_5_a_bits_mask),
		.auto_out_5_a_bits_data(out_xbar_auto_out_5_a_bits_data),
		.auto_out_5_d_ready(out_xbar_auto_out_5_d_ready),
		.auto_out_5_d_valid(out_xbar_auto_out_5_d_valid),
		.auto_out_5_d_bits_opcode(out_xbar_auto_out_5_d_bits_opcode),
		.auto_out_5_d_bits_param(out_xbar_auto_out_5_d_bits_param),
		.auto_out_5_d_bits_size(out_xbar_auto_out_5_d_bits_size),
		.auto_out_5_d_bits_source(out_xbar_auto_out_5_d_bits_source),
		.auto_out_5_d_bits_sink(out_xbar_auto_out_5_d_bits_sink),
		.auto_out_5_d_bits_denied(out_xbar_auto_out_5_d_bits_denied),
		.auto_out_5_d_bits_data(out_xbar_auto_out_5_d_bits_data),
		.auto_out_5_d_bits_corrupt(out_xbar_auto_out_5_d_bits_corrupt),
		.auto_out_4_a_ready(out_xbar_auto_out_4_a_ready),
		.auto_out_4_a_valid(out_xbar_auto_out_4_a_valid),
		.auto_out_4_a_bits_opcode(out_xbar_auto_out_4_a_bits_opcode),
		.auto_out_4_a_bits_param(out_xbar_auto_out_4_a_bits_param),
		.auto_out_4_a_bits_size(out_xbar_auto_out_4_a_bits_size),
		.auto_out_4_a_bits_source(out_xbar_auto_out_4_a_bits_source),
		.auto_out_4_a_bits_address(out_xbar_auto_out_4_a_bits_address),
		.auto_out_4_a_bits_mask(out_xbar_auto_out_4_a_bits_mask),
		.auto_out_4_a_bits_data(out_xbar_auto_out_4_a_bits_data),
		.auto_out_4_a_bits_corrupt(out_xbar_auto_out_4_a_bits_corrupt),
		.auto_out_4_d_ready(out_xbar_auto_out_4_d_ready),
		.auto_out_4_d_valid(out_xbar_auto_out_4_d_valid),
		.auto_out_4_d_bits_opcode(out_xbar_auto_out_4_d_bits_opcode),
		.auto_out_4_d_bits_size(out_xbar_auto_out_4_d_bits_size),
		.auto_out_4_d_bits_source(out_xbar_auto_out_4_d_bits_source),
		.auto_out_4_d_bits_data(out_xbar_auto_out_4_d_bits_data),
		.auto_out_3_a_ready(out_xbar_auto_out_3_a_ready),
		.auto_out_3_a_valid(out_xbar_auto_out_3_a_valid),
		.auto_out_3_a_bits_opcode(out_xbar_auto_out_3_a_bits_opcode),
		.auto_out_3_a_bits_param(out_xbar_auto_out_3_a_bits_param),
		.auto_out_3_a_bits_size(out_xbar_auto_out_3_a_bits_size),
		.auto_out_3_a_bits_source(out_xbar_auto_out_3_a_bits_source),
		.auto_out_3_a_bits_address(out_xbar_auto_out_3_a_bits_address),
		.auto_out_3_a_bits_mask(out_xbar_auto_out_3_a_bits_mask),
		.auto_out_3_a_bits_data(out_xbar_auto_out_3_a_bits_data),
		.auto_out_3_a_bits_corrupt(out_xbar_auto_out_3_a_bits_corrupt),
		.auto_out_3_d_ready(out_xbar_auto_out_3_d_ready),
		.auto_out_3_d_valid(out_xbar_auto_out_3_d_valid),
		.auto_out_3_d_bits_opcode(out_xbar_auto_out_3_d_bits_opcode),
		.auto_out_3_d_bits_size(out_xbar_auto_out_3_d_bits_size),
		.auto_out_3_d_bits_source(out_xbar_auto_out_3_d_bits_source),
		.auto_out_3_d_bits_data(out_xbar_auto_out_3_d_bits_data),
		.auto_out_2_a_ready(out_xbar_auto_out_2_a_ready),
		.auto_out_2_a_valid(out_xbar_auto_out_2_a_valid),
		.auto_out_2_a_bits_opcode(out_xbar_auto_out_2_a_bits_opcode),
		.auto_out_2_a_bits_param(out_xbar_auto_out_2_a_bits_param),
		.auto_out_2_a_bits_size(out_xbar_auto_out_2_a_bits_size),
		.auto_out_2_a_bits_source(out_xbar_auto_out_2_a_bits_source),
		.auto_out_2_a_bits_address(out_xbar_auto_out_2_a_bits_address),
		.auto_out_2_a_bits_mask(out_xbar_auto_out_2_a_bits_mask),
		.auto_out_2_a_bits_data(out_xbar_auto_out_2_a_bits_data),
		.auto_out_2_a_bits_corrupt(out_xbar_auto_out_2_a_bits_corrupt),
		.auto_out_2_d_ready(out_xbar_auto_out_2_d_ready),
		.auto_out_2_d_valid(out_xbar_auto_out_2_d_valid),
		.auto_out_2_d_bits_opcode(out_xbar_auto_out_2_d_bits_opcode),
		.auto_out_2_d_bits_size(out_xbar_auto_out_2_d_bits_size),
		.auto_out_2_d_bits_source(out_xbar_auto_out_2_d_bits_source),
		.auto_out_2_d_bits_data(out_xbar_auto_out_2_d_bits_data),
		.auto_out_1_a_ready(out_xbar_auto_out_1_a_ready),
		.auto_out_1_a_valid(out_xbar_auto_out_1_a_valid),
		.auto_out_1_a_bits_opcode(out_xbar_auto_out_1_a_bits_opcode),
		.auto_out_1_a_bits_param(out_xbar_auto_out_1_a_bits_param),
		.auto_out_1_a_bits_size(out_xbar_auto_out_1_a_bits_size),
		.auto_out_1_a_bits_source(out_xbar_auto_out_1_a_bits_source),
		.auto_out_1_a_bits_address(out_xbar_auto_out_1_a_bits_address),
		.auto_out_1_a_bits_mask(out_xbar_auto_out_1_a_bits_mask),
		.auto_out_1_a_bits_data(out_xbar_auto_out_1_a_bits_data),
		.auto_out_1_a_bits_corrupt(out_xbar_auto_out_1_a_bits_corrupt),
		.auto_out_1_d_ready(out_xbar_auto_out_1_d_ready),
		.auto_out_1_d_valid(out_xbar_auto_out_1_d_valid),
		.auto_out_1_d_bits_opcode(out_xbar_auto_out_1_d_bits_opcode),
		.auto_out_1_d_bits_param(out_xbar_auto_out_1_d_bits_param),
		.auto_out_1_d_bits_size(out_xbar_auto_out_1_d_bits_size),
		.auto_out_1_d_bits_source(out_xbar_auto_out_1_d_bits_source),
		.auto_out_1_d_bits_sink(out_xbar_auto_out_1_d_bits_sink),
		.auto_out_1_d_bits_denied(out_xbar_auto_out_1_d_bits_denied),
		.auto_out_1_d_bits_data(out_xbar_auto_out_1_d_bits_data),
		.auto_out_1_d_bits_corrupt(out_xbar_auto_out_1_d_bits_corrupt),
		.auto_out_0_a_ready(out_xbar_auto_out_0_a_ready),
		.auto_out_0_a_valid(out_xbar_auto_out_0_a_valid),
		.auto_out_0_a_bits_opcode(out_xbar_auto_out_0_a_bits_opcode),
		.auto_out_0_a_bits_param(out_xbar_auto_out_0_a_bits_param),
		.auto_out_0_a_bits_size(out_xbar_auto_out_0_a_bits_size),
		.auto_out_0_a_bits_source(out_xbar_auto_out_0_a_bits_source),
		.auto_out_0_a_bits_address(out_xbar_auto_out_0_a_bits_address),
		.auto_out_0_a_bits_mask(out_xbar_auto_out_0_a_bits_mask),
		.auto_out_0_a_bits_corrupt(out_xbar_auto_out_0_a_bits_corrupt),
		.auto_out_0_d_ready(out_xbar_auto_out_0_d_ready),
		.auto_out_0_d_valid(out_xbar_auto_out_0_d_valid),
		.auto_out_0_d_bits_opcode(out_xbar_auto_out_0_d_bits_opcode),
		.auto_out_0_d_bits_param(out_xbar_auto_out_0_d_bits_param),
		.auto_out_0_d_bits_size(out_xbar_auto_out_0_d_bits_size),
		.auto_out_0_d_bits_source(out_xbar_auto_out_0_d_bits_source),
		.auto_out_0_d_bits_sink(out_xbar_auto_out_0_d_bits_sink),
		.auto_out_0_d_bits_denied(out_xbar_auto_out_0_d_bits_denied),
		.auto_out_0_d_bits_data(out_xbar_auto_out_0_d_bits_data),
		.auto_out_0_d_bits_corrupt(out_xbar_auto_out_0_d_bits_corrupt)
	);
	TLBuffer_6 buffer(
		.clock(buffer_clock),
		.reset(buffer_reset),
		.auto_in_a_ready(buffer_auto_in_a_ready),
		.auto_in_a_valid(buffer_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_auto_in_d_ready),
		.auto_in_d_valid(buffer_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_auto_out_a_ready),
		.auto_out_a_valid(buffer_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_auto_out_d_ready),
		.auto_out_d_valid(buffer_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(buffer_auto_out_d_bits_param),
		.auto_out_d_bits_size(buffer_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_auto_out_d_bits_source),
		.auto_out_d_bits_sink(buffer_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
		.auto_out_d_bits_data(buffer_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt)
	);
	TLAtomicAutomata_1 atomics(
		.clock(atomics_clock),
		.reset(atomics_reset),
		.auto_in_a_ready(atomics_auto_in_a_ready),
		.auto_in_a_valid(atomics_auto_in_a_valid),
		.auto_in_a_bits_opcode(atomics_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(atomics_auto_in_a_bits_param),
		.auto_in_a_bits_size(atomics_auto_in_a_bits_size),
		.auto_in_a_bits_source(atomics_auto_in_a_bits_source),
		.auto_in_a_bits_address(atomics_auto_in_a_bits_address),
		.auto_in_a_bits_mask(atomics_auto_in_a_bits_mask),
		.auto_in_a_bits_data(atomics_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(atomics_auto_in_a_bits_corrupt),
		.auto_in_d_ready(atomics_auto_in_d_ready),
		.auto_in_d_valid(atomics_auto_in_d_valid),
		.auto_in_d_bits_opcode(atomics_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(atomics_auto_in_d_bits_param),
		.auto_in_d_bits_size(atomics_auto_in_d_bits_size),
		.auto_in_d_bits_source(atomics_auto_in_d_bits_source),
		.auto_in_d_bits_sink(atomics_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(atomics_auto_in_d_bits_denied),
		.auto_in_d_bits_data(atomics_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(atomics_auto_in_d_bits_corrupt),
		.auto_out_a_ready(atomics_auto_out_a_ready),
		.auto_out_a_valid(atomics_auto_out_a_valid),
		.auto_out_a_bits_opcode(atomics_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(atomics_auto_out_a_bits_param),
		.auto_out_a_bits_size(atomics_auto_out_a_bits_size),
		.auto_out_a_bits_source(atomics_auto_out_a_bits_source),
		.auto_out_a_bits_address(atomics_auto_out_a_bits_address),
		.auto_out_a_bits_mask(atomics_auto_out_a_bits_mask),
		.auto_out_a_bits_data(atomics_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(atomics_auto_out_a_bits_corrupt),
		.auto_out_d_ready(atomics_auto_out_d_ready),
		.auto_out_d_valid(atomics_auto_out_d_valid),
		.auto_out_d_bits_opcode(atomics_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(atomics_auto_out_d_bits_param),
		.auto_out_d_bits_size(atomics_auto_out_d_bits_size),
		.auto_out_d_bits_source(atomics_auto_out_d_bits_source),
		.auto_out_d_bits_sink(atomics_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(atomics_auto_out_d_bits_denied),
		.auto_out_d_bits_data(atomics_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(atomics_auto_out_d_bits_corrupt)
	);
	ErrorDeviceWrapper wrapped_error_device(
		.clock(wrapped_error_device_clock),
		.reset(wrapped_error_device_reset),
		.auto_buffer_in_a_ready(wrapped_error_device_auto_buffer_in_a_ready),
		.auto_buffer_in_a_valid(wrapped_error_device_auto_buffer_in_a_valid),
		.auto_buffer_in_a_bits_opcode(wrapped_error_device_auto_buffer_in_a_bits_opcode),
		.auto_buffer_in_a_bits_param(wrapped_error_device_auto_buffer_in_a_bits_param),
		.auto_buffer_in_a_bits_size(wrapped_error_device_auto_buffer_in_a_bits_size),
		.auto_buffer_in_a_bits_source(wrapped_error_device_auto_buffer_in_a_bits_source),
		.auto_buffer_in_a_bits_address(wrapped_error_device_auto_buffer_in_a_bits_address),
		.auto_buffer_in_a_bits_mask(wrapped_error_device_auto_buffer_in_a_bits_mask),
		.auto_buffer_in_a_bits_corrupt(wrapped_error_device_auto_buffer_in_a_bits_corrupt),
		.auto_buffer_in_d_ready(wrapped_error_device_auto_buffer_in_d_ready),
		.auto_buffer_in_d_valid(wrapped_error_device_auto_buffer_in_d_valid),
		.auto_buffer_in_d_bits_opcode(wrapped_error_device_auto_buffer_in_d_bits_opcode),
		.auto_buffer_in_d_bits_param(wrapped_error_device_auto_buffer_in_d_bits_param),
		.auto_buffer_in_d_bits_size(wrapped_error_device_auto_buffer_in_d_bits_size),
		.auto_buffer_in_d_bits_source(wrapped_error_device_auto_buffer_in_d_bits_source),
		.auto_buffer_in_d_bits_sink(wrapped_error_device_auto_buffer_in_d_bits_sink),
		.auto_buffer_in_d_bits_denied(wrapped_error_device_auto_buffer_in_d_bits_denied),
		.auto_buffer_in_d_bits_data(wrapped_error_device_auto_buffer_in_d_bits_data),
		.auto_buffer_in_d_bits_corrupt(wrapped_error_device_auto_buffer_in_d_bits_corrupt)
	);
	TLBuffer_8 buffer_1(
		.auto_in_a_ready(buffer_1_auto_in_a_ready),
		.auto_in_a_valid(buffer_1_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_1_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_1_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_1_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_1_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_1_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_1_auto_in_d_ready),
		.auto_in_d_valid(buffer_1_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_1_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_1_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_1_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_1_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_1_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_1_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_1_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_1_auto_out_a_ready),
		.auto_out_a_valid(buffer_1_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_1_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_1_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_1_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_1_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_1_auto_out_d_ready),
		.auto_out_d_valid(buffer_1_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(buffer_1_auto_out_d_bits_param),
		.auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
		.auto_out_d_bits_sink(buffer_1_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
		.auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt)
	);
	TLInterconnectCoupler_9 coupler_to_bus_named_subsystem_pbus(
		.auto_widget_in_a_ready(coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_ready),
		.auto_widget_in_a_valid(coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_valid),
		.auto_widget_in_a_bits_opcode(coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_opcode),
		.auto_widget_in_a_bits_param(coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_param),
		.auto_widget_in_a_bits_size(coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_size),
		.auto_widget_in_a_bits_source(coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_source),
		.auto_widget_in_a_bits_address(coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_address),
		.auto_widget_in_a_bits_mask(coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_mask),
		.auto_widget_in_a_bits_data(coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_data),
		.auto_widget_in_a_bits_corrupt(coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_corrupt),
		.auto_widget_in_d_ready(coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_ready),
		.auto_widget_in_d_valid(coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_valid),
		.auto_widget_in_d_bits_opcode(coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_opcode),
		.auto_widget_in_d_bits_param(coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_param),
		.auto_widget_in_d_bits_size(coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_size),
		.auto_widget_in_d_bits_source(coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_source),
		.auto_widget_in_d_bits_sink(coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_sink),
		.auto_widget_in_d_bits_denied(coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_denied),
		.auto_widget_in_d_bits_data(coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_data),
		.auto_widget_in_d_bits_corrupt(coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_corrupt),
		.auto_bus_xing_out_a_ready(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_ready),
		.auto_bus_xing_out_a_valid(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_valid),
		.auto_bus_xing_out_a_bits_opcode(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_opcode),
		.auto_bus_xing_out_a_bits_param(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_param),
		.auto_bus_xing_out_a_bits_size(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_size),
		.auto_bus_xing_out_a_bits_source(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_source),
		.auto_bus_xing_out_a_bits_address(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_address),
		.auto_bus_xing_out_a_bits_mask(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_mask),
		.auto_bus_xing_out_a_bits_data(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_data),
		.auto_bus_xing_out_a_bits_corrupt(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_corrupt),
		.auto_bus_xing_out_d_ready(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_ready),
		.auto_bus_xing_out_d_valid(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_valid),
		.auto_bus_xing_out_d_bits_opcode(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_opcode),
		.auto_bus_xing_out_d_bits_param(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_param),
		.auto_bus_xing_out_d_bits_size(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_size),
		.auto_bus_xing_out_d_bits_source(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_source),
		.auto_bus_xing_out_d_bits_sink(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_sink),
		.auto_bus_xing_out_d_bits_denied(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_denied),
		.auto_bus_xing_out_d_bits_data(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_data),
		.auto_bus_xing_out_d_bits_corrupt(coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_corrupt)
	);
	TLInterconnectCoupler_10 coupler_to_plic(
		.clock(coupler_to_plic_clock),
		.reset(coupler_to_plic_reset),
		.auto_fragmenter_out_a_ready(coupler_to_plic_auto_fragmenter_out_a_ready),
		.auto_fragmenter_out_a_valid(coupler_to_plic_auto_fragmenter_out_a_valid),
		.auto_fragmenter_out_a_bits_opcode(coupler_to_plic_auto_fragmenter_out_a_bits_opcode),
		.auto_fragmenter_out_a_bits_param(coupler_to_plic_auto_fragmenter_out_a_bits_param),
		.auto_fragmenter_out_a_bits_size(coupler_to_plic_auto_fragmenter_out_a_bits_size),
		.auto_fragmenter_out_a_bits_source(coupler_to_plic_auto_fragmenter_out_a_bits_source),
		.auto_fragmenter_out_a_bits_address(coupler_to_plic_auto_fragmenter_out_a_bits_address),
		.auto_fragmenter_out_a_bits_mask(coupler_to_plic_auto_fragmenter_out_a_bits_mask),
		.auto_fragmenter_out_a_bits_data(coupler_to_plic_auto_fragmenter_out_a_bits_data),
		.auto_fragmenter_out_a_bits_corrupt(coupler_to_plic_auto_fragmenter_out_a_bits_corrupt),
		.auto_fragmenter_out_d_ready(coupler_to_plic_auto_fragmenter_out_d_ready),
		.auto_fragmenter_out_d_valid(coupler_to_plic_auto_fragmenter_out_d_valid),
		.auto_fragmenter_out_d_bits_opcode(coupler_to_plic_auto_fragmenter_out_d_bits_opcode),
		.auto_fragmenter_out_d_bits_size(coupler_to_plic_auto_fragmenter_out_d_bits_size),
		.auto_fragmenter_out_d_bits_source(coupler_to_plic_auto_fragmenter_out_d_bits_source),
		.auto_fragmenter_out_d_bits_data(coupler_to_plic_auto_fragmenter_out_d_bits_data),
		.auto_tl_in_a_ready(coupler_to_plic_auto_tl_in_a_ready),
		.auto_tl_in_a_valid(coupler_to_plic_auto_tl_in_a_valid),
		.auto_tl_in_a_bits_opcode(coupler_to_plic_auto_tl_in_a_bits_opcode),
		.auto_tl_in_a_bits_param(coupler_to_plic_auto_tl_in_a_bits_param),
		.auto_tl_in_a_bits_size(coupler_to_plic_auto_tl_in_a_bits_size),
		.auto_tl_in_a_bits_source(coupler_to_plic_auto_tl_in_a_bits_source),
		.auto_tl_in_a_bits_address(coupler_to_plic_auto_tl_in_a_bits_address),
		.auto_tl_in_a_bits_mask(coupler_to_plic_auto_tl_in_a_bits_mask),
		.auto_tl_in_a_bits_data(coupler_to_plic_auto_tl_in_a_bits_data),
		.auto_tl_in_a_bits_corrupt(coupler_to_plic_auto_tl_in_a_bits_corrupt),
		.auto_tl_in_d_ready(coupler_to_plic_auto_tl_in_d_ready),
		.auto_tl_in_d_valid(coupler_to_plic_auto_tl_in_d_valid),
		.auto_tl_in_d_bits_opcode(coupler_to_plic_auto_tl_in_d_bits_opcode),
		.auto_tl_in_d_bits_size(coupler_to_plic_auto_tl_in_d_bits_size),
		.auto_tl_in_d_bits_source(coupler_to_plic_auto_tl_in_d_bits_source),
		.auto_tl_in_d_bits_data(coupler_to_plic_auto_tl_in_d_bits_data)
	);
	TLInterconnectCoupler_11 coupler_to_clint(
		.clock(coupler_to_clint_clock),
		.reset(coupler_to_clint_reset),
		.auto_fragmenter_out_a_ready(coupler_to_clint_auto_fragmenter_out_a_ready),
		.auto_fragmenter_out_a_valid(coupler_to_clint_auto_fragmenter_out_a_valid),
		.auto_fragmenter_out_a_bits_opcode(coupler_to_clint_auto_fragmenter_out_a_bits_opcode),
		.auto_fragmenter_out_a_bits_param(coupler_to_clint_auto_fragmenter_out_a_bits_param),
		.auto_fragmenter_out_a_bits_size(coupler_to_clint_auto_fragmenter_out_a_bits_size),
		.auto_fragmenter_out_a_bits_source(coupler_to_clint_auto_fragmenter_out_a_bits_source),
		.auto_fragmenter_out_a_bits_address(coupler_to_clint_auto_fragmenter_out_a_bits_address),
		.auto_fragmenter_out_a_bits_mask(coupler_to_clint_auto_fragmenter_out_a_bits_mask),
		.auto_fragmenter_out_a_bits_data(coupler_to_clint_auto_fragmenter_out_a_bits_data),
		.auto_fragmenter_out_a_bits_corrupt(coupler_to_clint_auto_fragmenter_out_a_bits_corrupt),
		.auto_fragmenter_out_d_ready(coupler_to_clint_auto_fragmenter_out_d_ready),
		.auto_fragmenter_out_d_valid(coupler_to_clint_auto_fragmenter_out_d_valid),
		.auto_fragmenter_out_d_bits_opcode(coupler_to_clint_auto_fragmenter_out_d_bits_opcode),
		.auto_fragmenter_out_d_bits_size(coupler_to_clint_auto_fragmenter_out_d_bits_size),
		.auto_fragmenter_out_d_bits_source(coupler_to_clint_auto_fragmenter_out_d_bits_source),
		.auto_fragmenter_out_d_bits_data(coupler_to_clint_auto_fragmenter_out_d_bits_data),
		.auto_tl_in_a_ready(coupler_to_clint_auto_tl_in_a_ready),
		.auto_tl_in_a_valid(coupler_to_clint_auto_tl_in_a_valid),
		.auto_tl_in_a_bits_opcode(coupler_to_clint_auto_tl_in_a_bits_opcode),
		.auto_tl_in_a_bits_param(coupler_to_clint_auto_tl_in_a_bits_param),
		.auto_tl_in_a_bits_size(coupler_to_clint_auto_tl_in_a_bits_size),
		.auto_tl_in_a_bits_source(coupler_to_clint_auto_tl_in_a_bits_source),
		.auto_tl_in_a_bits_address(coupler_to_clint_auto_tl_in_a_bits_address),
		.auto_tl_in_a_bits_mask(coupler_to_clint_auto_tl_in_a_bits_mask),
		.auto_tl_in_a_bits_data(coupler_to_clint_auto_tl_in_a_bits_data),
		.auto_tl_in_a_bits_corrupt(coupler_to_clint_auto_tl_in_a_bits_corrupt),
		.auto_tl_in_d_ready(coupler_to_clint_auto_tl_in_d_ready),
		.auto_tl_in_d_valid(coupler_to_clint_auto_tl_in_d_valid),
		.auto_tl_in_d_bits_opcode(coupler_to_clint_auto_tl_in_d_bits_opcode),
		.auto_tl_in_d_bits_size(coupler_to_clint_auto_tl_in_d_bits_size),
		.auto_tl_in_d_bits_source(coupler_to_clint_auto_tl_in_d_bits_source),
		.auto_tl_in_d_bits_data(coupler_to_clint_auto_tl_in_d_bits_data)
	);
	TLInterconnectCoupler_12 coupler_to_debug(
		.clock(coupler_to_debug_clock),
		.reset(coupler_to_debug_reset),
		.auto_fragmenter_out_a_ready(coupler_to_debug_auto_fragmenter_out_a_ready),
		.auto_fragmenter_out_a_valid(coupler_to_debug_auto_fragmenter_out_a_valid),
		.auto_fragmenter_out_a_bits_opcode(coupler_to_debug_auto_fragmenter_out_a_bits_opcode),
		.auto_fragmenter_out_a_bits_param(coupler_to_debug_auto_fragmenter_out_a_bits_param),
		.auto_fragmenter_out_a_bits_size(coupler_to_debug_auto_fragmenter_out_a_bits_size),
		.auto_fragmenter_out_a_bits_source(coupler_to_debug_auto_fragmenter_out_a_bits_source),
		.auto_fragmenter_out_a_bits_address(coupler_to_debug_auto_fragmenter_out_a_bits_address),
		.auto_fragmenter_out_a_bits_mask(coupler_to_debug_auto_fragmenter_out_a_bits_mask),
		.auto_fragmenter_out_a_bits_data(coupler_to_debug_auto_fragmenter_out_a_bits_data),
		.auto_fragmenter_out_a_bits_corrupt(coupler_to_debug_auto_fragmenter_out_a_bits_corrupt),
		.auto_fragmenter_out_d_ready(coupler_to_debug_auto_fragmenter_out_d_ready),
		.auto_fragmenter_out_d_valid(coupler_to_debug_auto_fragmenter_out_d_valid),
		.auto_fragmenter_out_d_bits_opcode(coupler_to_debug_auto_fragmenter_out_d_bits_opcode),
		.auto_fragmenter_out_d_bits_size(coupler_to_debug_auto_fragmenter_out_d_bits_size),
		.auto_fragmenter_out_d_bits_source(coupler_to_debug_auto_fragmenter_out_d_bits_source),
		.auto_fragmenter_out_d_bits_data(coupler_to_debug_auto_fragmenter_out_d_bits_data),
		.auto_tl_in_a_ready(coupler_to_debug_auto_tl_in_a_ready),
		.auto_tl_in_a_valid(coupler_to_debug_auto_tl_in_a_valid),
		.auto_tl_in_a_bits_opcode(coupler_to_debug_auto_tl_in_a_bits_opcode),
		.auto_tl_in_a_bits_param(coupler_to_debug_auto_tl_in_a_bits_param),
		.auto_tl_in_a_bits_size(coupler_to_debug_auto_tl_in_a_bits_size),
		.auto_tl_in_a_bits_source(coupler_to_debug_auto_tl_in_a_bits_source),
		.auto_tl_in_a_bits_address(coupler_to_debug_auto_tl_in_a_bits_address),
		.auto_tl_in_a_bits_mask(coupler_to_debug_auto_tl_in_a_bits_mask),
		.auto_tl_in_a_bits_data(coupler_to_debug_auto_tl_in_a_bits_data),
		.auto_tl_in_a_bits_corrupt(coupler_to_debug_auto_tl_in_a_bits_corrupt),
		.auto_tl_in_d_ready(coupler_to_debug_auto_tl_in_d_ready),
		.auto_tl_in_d_valid(coupler_to_debug_auto_tl_in_d_valid),
		.auto_tl_in_d_bits_opcode(coupler_to_debug_auto_tl_in_d_bits_opcode),
		.auto_tl_in_d_bits_size(coupler_to_debug_auto_tl_in_d_bits_size),
		.auto_tl_in_d_bits_source(coupler_to_debug_auto_tl_in_d_bits_source),
		.auto_tl_in_d_bits_data(coupler_to_debug_auto_tl_in_d_bits_data)
	);
	TLInterconnectCoupler_13 coupler_to_tile(
		.auto_tl_slave_clock_xing_out_a_ready(coupler_to_tile_auto_tl_slave_clock_xing_out_a_ready),
		.auto_tl_slave_clock_xing_out_a_valid(coupler_to_tile_auto_tl_slave_clock_xing_out_a_valid),
		.auto_tl_slave_clock_xing_out_a_bits_opcode(coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_opcode),
		.auto_tl_slave_clock_xing_out_a_bits_param(coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_param),
		.auto_tl_slave_clock_xing_out_a_bits_size(coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_size),
		.auto_tl_slave_clock_xing_out_a_bits_source(coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_source),
		.auto_tl_slave_clock_xing_out_a_bits_address(coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_address),
		.auto_tl_slave_clock_xing_out_a_bits_mask(coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_mask),
		.auto_tl_slave_clock_xing_out_a_bits_data(coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_data),
		.auto_tl_slave_clock_xing_out_d_ready(coupler_to_tile_auto_tl_slave_clock_xing_out_d_ready),
		.auto_tl_slave_clock_xing_out_d_valid(coupler_to_tile_auto_tl_slave_clock_xing_out_d_valid),
		.auto_tl_slave_clock_xing_out_d_bits_opcode(coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_opcode),
		.auto_tl_slave_clock_xing_out_d_bits_param(coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_param),
		.auto_tl_slave_clock_xing_out_d_bits_size(coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_size),
		.auto_tl_slave_clock_xing_out_d_bits_source(coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_source),
		.auto_tl_slave_clock_xing_out_d_bits_sink(coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_sink),
		.auto_tl_slave_clock_xing_out_d_bits_denied(coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_denied),
		.auto_tl_slave_clock_xing_out_d_bits_data(coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_data),
		.auto_tl_slave_clock_xing_out_d_bits_corrupt(coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_corrupt),
		.auto_tl_in_a_ready(coupler_to_tile_auto_tl_in_a_ready),
		.auto_tl_in_a_valid(coupler_to_tile_auto_tl_in_a_valid),
		.auto_tl_in_a_bits_opcode(coupler_to_tile_auto_tl_in_a_bits_opcode),
		.auto_tl_in_a_bits_param(coupler_to_tile_auto_tl_in_a_bits_param),
		.auto_tl_in_a_bits_size(coupler_to_tile_auto_tl_in_a_bits_size),
		.auto_tl_in_a_bits_source(coupler_to_tile_auto_tl_in_a_bits_source),
		.auto_tl_in_a_bits_address(coupler_to_tile_auto_tl_in_a_bits_address),
		.auto_tl_in_a_bits_mask(coupler_to_tile_auto_tl_in_a_bits_mask),
		.auto_tl_in_a_bits_data(coupler_to_tile_auto_tl_in_a_bits_data),
		.auto_tl_in_d_ready(coupler_to_tile_auto_tl_in_d_ready),
		.auto_tl_in_d_valid(coupler_to_tile_auto_tl_in_d_valid),
		.auto_tl_in_d_bits_opcode(coupler_to_tile_auto_tl_in_d_bits_opcode),
		.auto_tl_in_d_bits_param(coupler_to_tile_auto_tl_in_d_bits_param),
		.auto_tl_in_d_bits_size(coupler_to_tile_auto_tl_in_d_bits_size),
		.auto_tl_in_d_bits_source(coupler_to_tile_auto_tl_in_d_bits_source),
		.auto_tl_in_d_bits_sink(coupler_to_tile_auto_tl_in_d_bits_sink),
		.auto_tl_in_d_bits_denied(coupler_to_tile_auto_tl_in_d_bits_denied),
		.auto_tl_in_d_bits_data(coupler_to_tile_auto_tl_in_d_bits_data),
		.auto_tl_in_d_bits_corrupt(coupler_to_tile_auto_tl_in_d_bits_corrupt)
	);
	TLInterconnectCoupler_14 coupler_to_bootrom(
		.clock(coupler_to_bootrom_clock),
		.reset(coupler_to_bootrom_reset),
		.auto_fragmenter_out_a_ready(coupler_to_bootrom_auto_fragmenter_out_a_ready),
		.auto_fragmenter_out_a_valid(coupler_to_bootrom_auto_fragmenter_out_a_valid),
		.auto_fragmenter_out_a_bits_opcode(coupler_to_bootrom_auto_fragmenter_out_a_bits_opcode),
		.auto_fragmenter_out_a_bits_param(coupler_to_bootrom_auto_fragmenter_out_a_bits_param),
		.auto_fragmenter_out_a_bits_size(coupler_to_bootrom_auto_fragmenter_out_a_bits_size),
		.auto_fragmenter_out_a_bits_source(coupler_to_bootrom_auto_fragmenter_out_a_bits_source),
		.auto_fragmenter_out_a_bits_address(coupler_to_bootrom_auto_fragmenter_out_a_bits_address),
		.auto_fragmenter_out_a_bits_mask(coupler_to_bootrom_auto_fragmenter_out_a_bits_mask),
		.auto_fragmenter_out_a_bits_corrupt(coupler_to_bootrom_auto_fragmenter_out_a_bits_corrupt),
		.auto_fragmenter_out_d_ready(coupler_to_bootrom_auto_fragmenter_out_d_ready),
		.auto_fragmenter_out_d_valid(coupler_to_bootrom_auto_fragmenter_out_d_valid),
		.auto_fragmenter_out_d_bits_size(coupler_to_bootrom_auto_fragmenter_out_d_bits_size),
		.auto_fragmenter_out_d_bits_source(coupler_to_bootrom_auto_fragmenter_out_d_bits_source),
		.auto_fragmenter_out_d_bits_data(coupler_to_bootrom_auto_fragmenter_out_d_bits_data),
		.auto_tl_in_a_ready(coupler_to_bootrom_auto_tl_in_a_ready),
		.auto_tl_in_a_valid(coupler_to_bootrom_auto_tl_in_a_valid),
		.auto_tl_in_a_bits_opcode(coupler_to_bootrom_auto_tl_in_a_bits_opcode),
		.auto_tl_in_a_bits_param(coupler_to_bootrom_auto_tl_in_a_bits_param),
		.auto_tl_in_a_bits_size(coupler_to_bootrom_auto_tl_in_a_bits_size),
		.auto_tl_in_a_bits_source(coupler_to_bootrom_auto_tl_in_a_bits_source),
		.auto_tl_in_a_bits_address(coupler_to_bootrom_auto_tl_in_a_bits_address),
		.auto_tl_in_a_bits_mask(coupler_to_bootrom_auto_tl_in_a_bits_mask),
		.auto_tl_in_a_bits_corrupt(coupler_to_bootrom_auto_tl_in_a_bits_corrupt),
		.auto_tl_in_d_ready(coupler_to_bootrom_auto_tl_in_d_ready),
		.auto_tl_in_d_valid(coupler_to_bootrom_auto_tl_in_d_valid),
		.auto_tl_in_d_bits_size(coupler_to_bootrom_auto_tl_in_d_bits_size),
		.auto_tl_in_d_bits_source(coupler_to_bootrom_auto_tl_in_d_bits_source),
		.auto_tl_in_d_bits_data(coupler_to_bootrom_auto_tl_in_d_bits_data)
	);
	TLInterconnectCoupler_15 coupler_from_port_named_custom_boot_pin(
		.auto_tl_in_a_ready(coupler_from_port_named_custom_boot_pin_auto_tl_in_a_ready),
		.auto_tl_in_a_valid(coupler_from_port_named_custom_boot_pin_auto_tl_in_a_valid),
		.auto_tl_in_a_bits_address(coupler_from_port_named_custom_boot_pin_auto_tl_in_a_bits_address),
		.auto_tl_in_a_bits_data(coupler_from_port_named_custom_boot_pin_auto_tl_in_a_bits_data),
		.auto_tl_in_d_valid(coupler_from_port_named_custom_boot_pin_auto_tl_in_d_valid),
		.auto_tl_out_a_ready(coupler_from_port_named_custom_boot_pin_auto_tl_out_a_ready),
		.auto_tl_out_a_valid(coupler_from_port_named_custom_boot_pin_auto_tl_out_a_valid),
		.auto_tl_out_a_bits_address(coupler_from_port_named_custom_boot_pin_auto_tl_out_a_bits_address),
		.auto_tl_out_a_bits_data(coupler_from_port_named_custom_boot_pin_auto_tl_out_a_bits_data),
		.auto_tl_out_d_valid(coupler_from_port_named_custom_boot_pin_auto_tl_out_d_valid)
	);
	TLInterconnectCoupler_16 coupler_to_slave_named_clockgater(
		.clock(coupler_to_slave_named_clockgater_clock),
		.reset(coupler_to_slave_named_clockgater_reset),
		.auto_buffer_in_a_ready(coupler_to_slave_named_clockgater_auto_buffer_in_a_ready),
		.auto_buffer_in_a_valid(coupler_to_slave_named_clockgater_auto_buffer_in_a_valid),
		.auto_buffer_in_a_bits_opcode(coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_opcode),
		.auto_buffer_in_a_bits_param(coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_param),
		.auto_buffer_in_a_bits_size(coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_size),
		.auto_buffer_in_a_bits_source(coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_source),
		.auto_buffer_in_a_bits_address(coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_address),
		.auto_buffer_in_a_bits_mask(coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_mask),
		.auto_buffer_in_a_bits_data(coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_data),
		.auto_buffer_in_a_bits_corrupt(coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_corrupt),
		.auto_buffer_in_d_ready(coupler_to_slave_named_clockgater_auto_buffer_in_d_ready),
		.auto_buffer_in_d_valid(coupler_to_slave_named_clockgater_auto_buffer_in_d_valid),
		.auto_buffer_in_d_bits_opcode(coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_opcode),
		.auto_buffer_in_d_bits_param(coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_param),
		.auto_buffer_in_d_bits_size(coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_size),
		.auto_buffer_in_d_bits_source(coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_source),
		.auto_buffer_in_d_bits_sink(coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_sink),
		.auto_buffer_in_d_bits_denied(coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_denied),
		.auto_buffer_in_d_bits_data(coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_data),
		.auto_buffer_in_d_bits_corrupt(coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_corrupt),
		.auto_buffer_out_a_ready(coupler_to_slave_named_clockgater_auto_buffer_out_a_ready),
		.auto_buffer_out_a_valid(coupler_to_slave_named_clockgater_auto_buffer_out_a_valid),
		.auto_buffer_out_a_bits_opcode(coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_opcode),
		.auto_buffer_out_a_bits_param(coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_param),
		.auto_buffer_out_a_bits_size(coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_size),
		.auto_buffer_out_a_bits_source(coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_source),
		.auto_buffer_out_a_bits_address(coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_address),
		.auto_buffer_out_a_bits_mask(coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_mask),
		.auto_buffer_out_a_bits_data(coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_data),
		.auto_buffer_out_a_bits_corrupt(coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_corrupt),
		.auto_buffer_out_d_ready(coupler_to_slave_named_clockgater_auto_buffer_out_d_ready),
		.auto_buffer_out_d_valid(coupler_to_slave_named_clockgater_auto_buffer_out_d_valid),
		.auto_buffer_out_d_bits_opcode(coupler_to_slave_named_clockgater_auto_buffer_out_d_bits_opcode),
		.auto_buffer_out_d_bits_size(coupler_to_slave_named_clockgater_auto_buffer_out_d_bits_size),
		.auto_buffer_out_d_bits_source(coupler_to_slave_named_clockgater_auto_buffer_out_d_bits_source),
		.auto_buffer_out_d_bits_data(coupler_to_slave_named_clockgater_auto_buffer_out_d_bits_data)
	);
	TLInterconnectCoupler_17 coupler_to_slave_named_tileresetsetter(
		.clock(coupler_to_slave_named_tileresetsetter_clock),
		.reset(coupler_to_slave_named_tileresetsetter_reset),
		.auto_buffer_in_a_ready(coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_ready),
		.auto_buffer_in_a_valid(coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_valid),
		.auto_buffer_in_a_bits_opcode(coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_opcode),
		.auto_buffer_in_a_bits_param(coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_param),
		.auto_buffer_in_a_bits_size(coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_size),
		.auto_buffer_in_a_bits_source(coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_source),
		.auto_buffer_in_a_bits_address(coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_address),
		.auto_buffer_in_a_bits_mask(coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_mask),
		.auto_buffer_in_a_bits_data(coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_data),
		.auto_buffer_in_a_bits_corrupt(coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_corrupt),
		.auto_buffer_in_d_ready(coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_ready),
		.auto_buffer_in_d_valid(coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_valid),
		.auto_buffer_in_d_bits_opcode(coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_opcode),
		.auto_buffer_in_d_bits_param(coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_param),
		.auto_buffer_in_d_bits_size(coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_size),
		.auto_buffer_in_d_bits_source(coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_source),
		.auto_buffer_in_d_bits_sink(coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_sink),
		.auto_buffer_in_d_bits_denied(coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_denied),
		.auto_buffer_in_d_bits_data(coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_data),
		.auto_buffer_in_d_bits_corrupt(coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_corrupt),
		.auto_buffer_out_a_ready(coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_ready),
		.auto_buffer_out_a_valid(coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_valid),
		.auto_buffer_out_a_bits_opcode(coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_opcode),
		.auto_buffer_out_a_bits_param(coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_param),
		.auto_buffer_out_a_bits_size(coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_size),
		.auto_buffer_out_a_bits_source(coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_source),
		.auto_buffer_out_a_bits_address(coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_address),
		.auto_buffer_out_a_bits_mask(coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_mask),
		.auto_buffer_out_a_bits_data(coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_data),
		.auto_buffer_out_a_bits_corrupt(coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_corrupt),
		.auto_buffer_out_d_ready(coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_ready),
		.auto_buffer_out_d_valid(coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_valid),
		.auto_buffer_out_d_bits_opcode(coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_bits_opcode),
		.auto_buffer_out_d_bits_size(coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_bits_size),
		.auto_buffer_out_d_bits_source(coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_bits_source),
		.auto_buffer_out_d_bits_data(coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_bits_data)
	);
	assign auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_valid = coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_valid;
	assign auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_opcode = coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_opcode;
	assign auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_param = coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_param;
	assign auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_size = coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_size;
	assign auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_source = coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_source;
	assign auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_address = coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_address;
	assign auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_mask = coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_mask;
	assign auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_data = coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_data;
	assign auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_corrupt = coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_bits_corrupt;
	assign auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_ready = coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_ready;
	assign auto_coupler_to_slave_named_clockgater_buffer_out_a_valid = coupler_to_slave_named_clockgater_auto_buffer_out_a_valid;
	assign auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_opcode = coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_opcode;
	assign auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_param = coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_param;
	assign auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_size = coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_size;
	assign auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_source = coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_source;
	assign auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_address = coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_address;
	assign auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_mask = coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_mask;
	assign auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_data = coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_data;
	assign auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_corrupt = coupler_to_slave_named_clockgater_auto_buffer_out_a_bits_corrupt;
	assign auto_coupler_to_slave_named_clockgater_buffer_out_d_ready = coupler_to_slave_named_clockgater_auto_buffer_out_d_ready;
	assign auto_coupler_to_bootrom_fragmenter_out_a_valid = coupler_to_bootrom_auto_fragmenter_out_a_valid;
	assign auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode = coupler_to_bootrom_auto_fragmenter_out_a_bits_opcode;
	assign auto_coupler_to_bootrom_fragmenter_out_a_bits_param = coupler_to_bootrom_auto_fragmenter_out_a_bits_param;
	assign auto_coupler_to_bootrom_fragmenter_out_a_bits_size = coupler_to_bootrom_auto_fragmenter_out_a_bits_size;
	assign auto_coupler_to_bootrom_fragmenter_out_a_bits_source = coupler_to_bootrom_auto_fragmenter_out_a_bits_source;
	assign auto_coupler_to_bootrom_fragmenter_out_a_bits_address = coupler_to_bootrom_auto_fragmenter_out_a_bits_address;
	assign auto_coupler_to_bootrom_fragmenter_out_a_bits_mask = coupler_to_bootrom_auto_fragmenter_out_a_bits_mask;
	assign auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt = coupler_to_bootrom_auto_fragmenter_out_a_bits_corrupt;
	assign auto_coupler_to_bootrom_fragmenter_out_d_ready = coupler_to_bootrom_auto_fragmenter_out_d_ready;
	assign auto_coupler_to_tile_tl_slave_clock_xing_out_a_valid = coupler_to_tile_auto_tl_slave_clock_xing_out_a_valid;
	assign auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_opcode = coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_opcode;
	assign auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_param = coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_param;
	assign auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_size = coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_size;
	assign auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_source = coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_source;
	assign auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_address = coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_address;
	assign auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_mask = coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_mask;
	assign auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_data = coupler_to_tile_auto_tl_slave_clock_xing_out_a_bits_data;
	assign auto_coupler_to_tile_tl_slave_clock_xing_out_d_ready = coupler_to_tile_auto_tl_slave_clock_xing_out_d_ready;
	assign auto_coupler_to_debug_fragmenter_out_a_valid = coupler_to_debug_auto_fragmenter_out_a_valid;
	assign auto_coupler_to_debug_fragmenter_out_a_bits_opcode = coupler_to_debug_auto_fragmenter_out_a_bits_opcode;
	assign auto_coupler_to_debug_fragmenter_out_a_bits_param = coupler_to_debug_auto_fragmenter_out_a_bits_param;
	assign auto_coupler_to_debug_fragmenter_out_a_bits_size = coupler_to_debug_auto_fragmenter_out_a_bits_size;
	assign auto_coupler_to_debug_fragmenter_out_a_bits_source = coupler_to_debug_auto_fragmenter_out_a_bits_source;
	assign auto_coupler_to_debug_fragmenter_out_a_bits_address = coupler_to_debug_auto_fragmenter_out_a_bits_address;
	assign auto_coupler_to_debug_fragmenter_out_a_bits_mask = coupler_to_debug_auto_fragmenter_out_a_bits_mask;
	assign auto_coupler_to_debug_fragmenter_out_a_bits_data = coupler_to_debug_auto_fragmenter_out_a_bits_data;
	assign auto_coupler_to_debug_fragmenter_out_a_bits_corrupt = coupler_to_debug_auto_fragmenter_out_a_bits_corrupt;
	assign auto_coupler_to_debug_fragmenter_out_d_ready = coupler_to_debug_auto_fragmenter_out_d_ready;
	assign auto_coupler_to_clint_fragmenter_out_a_valid = coupler_to_clint_auto_fragmenter_out_a_valid;
	assign auto_coupler_to_clint_fragmenter_out_a_bits_opcode = coupler_to_clint_auto_fragmenter_out_a_bits_opcode;
	assign auto_coupler_to_clint_fragmenter_out_a_bits_param = coupler_to_clint_auto_fragmenter_out_a_bits_param;
	assign auto_coupler_to_clint_fragmenter_out_a_bits_size = coupler_to_clint_auto_fragmenter_out_a_bits_size;
	assign auto_coupler_to_clint_fragmenter_out_a_bits_source = coupler_to_clint_auto_fragmenter_out_a_bits_source;
	assign auto_coupler_to_clint_fragmenter_out_a_bits_address = coupler_to_clint_auto_fragmenter_out_a_bits_address;
	assign auto_coupler_to_clint_fragmenter_out_a_bits_mask = coupler_to_clint_auto_fragmenter_out_a_bits_mask;
	assign auto_coupler_to_clint_fragmenter_out_a_bits_data = coupler_to_clint_auto_fragmenter_out_a_bits_data;
	assign auto_coupler_to_clint_fragmenter_out_a_bits_corrupt = coupler_to_clint_auto_fragmenter_out_a_bits_corrupt;
	assign auto_coupler_to_clint_fragmenter_out_d_ready = coupler_to_clint_auto_fragmenter_out_d_ready;
	assign auto_coupler_to_plic_fragmenter_out_a_valid = coupler_to_plic_auto_fragmenter_out_a_valid;
	assign auto_coupler_to_plic_fragmenter_out_a_bits_opcode = coupler_to_plic_auto_fragmenter_out_a_bits_opcode;
	assign auto_coupler_to_plic_fragmenter_out_a_bits_param = coupler_to_plic_auto_fragmenter_out_a_bits_param;
	assign auto_coupler_to_plic_fragmenter_out_a_bits_size = coupler_to_plic_auto_fragmenter_out_a_bits_size;
	assign auto_coupler_to_plic_fragmenter_out_a_bits_source = coupler_to_plic_auto_fragmenter_out_a_bits_source;
	assign auto_coupler_to_plic_fragmenter_out_a_bits_address = coupler_to_plic_auto_fragmenter_out_a_bits_address;
	assign auto_coupler_to_plic_fragmenter_out_a_bits_mask = coupler_to_plic_auto_fragmenter_out_a_bits_mask;
	assign auto_coupler_to_plic_fragmenter_out_a_bits_data = coupler_to_plic_auto_fragmenter_out_a_bits_data;
	assign auto_coupler_to_plic_fragmenter_out_a_bits_corrupt = coupler_to_plic_auto_fragmenter_out_a_bits_corrupt;
	assign auto_coupler_to_plic_fragmenter_out_d_ready = coupler_to_plic_auto_fragmenter_out_d_ready;
	assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid = coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_valid;
	assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode = coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_opcode;
	assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param = coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_param;
	assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size = coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_size;
	assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source = coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_source;
	assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address = coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_address;
	assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask = coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_mask;
	assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data = coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_data;
	assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_corrupt = coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_corrupt;
	assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready = coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_ready;
	assign auto_fixedClockNode_out_4_clock = fixedClockNode_auto_out_5_clock;
	assign auto_fixedClockNode_out_4_reset = fixedClockNode_auto_out_5_reset;
	assign auto_fixedClockNode_out_3_clock = fixedClockNode_auto_out_4_clock;
	assign auto_fixedClockNode_out_3_reset = fixedClockNode_auto_out_4_reset;
	assign auto_fixedClockNode_out_2_clock = fixedClockNode_auto_out_3_clock;
	assign auto_fixedClockNode_out_2_reset = fixedClockNode_auto_out_3_reset;
	assign auto_fixedClockNode_out_0_clock = fixedClockNode_auto_out_1_clock;
	assign auto_fixedClockNode_out_0_reset = fixedClockNode_auto_out_1_reset;
	assign auto_bus_xing_in_a_ready = buffer_1_auto_in_a_ready;
	assign auto_bus_xing_in_d_valid = buffer_1_auto_in_d_valid;
	assign auto_bus_xing_in_d_bits_opcode = buffer_1_auto_in_d_bits_opcode;
	assign auto_bus_xing_in_d_bits_param = buffer_1_auto_in_d_bits_param;
	assign auto_bus_xing_in_d_bits_size = buffer_1_auto_in_d_bits_size;
	assign auto_bus_xing_in_d_bits_source = buffer_1_auto_in_d_bits_source;
	assign auto_bus_xing_in_d_bits_sink = buffer_1_auto_in_d_bits_sink;
	assign auto_bus_xing_in_d_bits_denied = buffer_1_auto_in_d_bits_denied;
	assign auto_bus_xing_in_d_bits_data = buffer_1_auto_in_d_bits_data;
	assign auto_bus_xing_in_d_bits_corrupt = buffer_1_auto_in_d_bits_corrupt;
	assign clock = fixedClockNode_auto_out_0_clock;
	assign reset = fixedClockNode_auto_out_0_reset;
	assign subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_clock = auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock;
	assign subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_reset = auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset;
	assign clockGroup_auto_in_member_subsystem_cbus_0_clock = subsystem_cbus_clock_groups_auto_out_member_subsystem_cbus_0_clock;
	assign clockGroup_auto_in_member_subsystem_cbus_0_reset = subsystem_cbus_clock_groups_auto_out_member_subsystem_cbus_0_reset;
	assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock;
	assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset;
	assign fixer_clock = fixedClockNode_auto_out_0_clock;
	assign fixer_reset = fixedClockNode_auto_out_0_reset;
	assign fixer_auto_in_a_valid = buffer_auto_out_a_valid;
	assign fixer_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode;
	assign fixer_auto_in_a_bits_param = buffer_auto_out_a_bits_param;
	assign fixer_auto_in_a_bits_size = buffer_auto_out_a_bits_size;
	assign fixer_auto_in_a_bits_source = buffer_auto_out_a_bits_source;
	assign fixer_auto_in_a_bits_address = buffer_auto_out_a_bits_address;
	assign fixer_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask;
	assign fixer_auto_in_a_bits_data = buffer_auto_out_a_bits_data;
	assign fixer_auto_in_a_bits_corrupt = buffer_auto_out_a_bits_corrupt;
	assign fixer_auto_in_d_ready = buffer_auto_out_d_ready;
	assign fixer_auto_out_a_ready = out_xbar_auto_in_a_ready;
	assign fixer_auto_out_d_valid = out_xbar_auto_in_d_valid;
	assign fixer_auto_out_d_bits_opcode = out_xbar_auto_in_d_bits_opcode;
	assign fixer_auto_out_d_bits_param = out_xbar_auto_in_d_bits_param;
	assign fixer_auto_out_d_bits_size = out_xbar_auto_in_d_bits_size;
	assign fixer_auto_out_d_bits_source = out_xbar_auto_in_d_bits_source;
	assign fixer_auto_out_d_bits_sink = out_xbar_auto_in_d_bits_sink;
	assign fixer_auto_out_d_bits_denied = out_xbar_auto_in_d_bits_denied;
	assign fixer_auto_out_d_bits_data = out_xbar_auto_in_d_bits_data;
	assign fixer_auto_out_d_bits_corrupt = out_xbar_auto_in_d_bits_corrupt;
	assign in_xbar_clock = fixedClockNode_auto_out_0_clock;
	assign in_xbar_reset = fixedClockNode_auto_out_0_reset;
	assign in_xbar_auto_in_1_a_valid = coupler_from_port_named_custom_boot_pin_auto_tl_out_a_valid;
	assign in_xbar_auto_in_1_a_bits_address = coupler_from_port_named_custom_boot_pin_auto_tl_out_a_bits_address;
	assign in_xbar_auto_in_1_a_bits_data = coupler_from_port_named_custom_boot_pin_auto_tl_out_a_bits_data;
	assign in_xbar_auto_in_0_a_valid = buffer_1_auto_out_a_valid;
	assign in_xbar_auto_in_0_a_bits_opcode = buffer_1_auto_out_a_bits_opcode;
	assign in_xbar_auto_in_0_a_bits_param = buffer_1_auto_out_a_bits_param;
	assign in_xbar_auto_in_0_a_bits_size = buffer_1_auto_out_a_bits_size;
	assign in_xbar_auto_in_0_a_bits_source = buffer_1_auto_out_a_bits_source;
	assign in_xbar_auto_in_0_a_bits_address = buffer_1_auto_out_a_bits_address;
	assign in_xbar_auto_in_0_a_bits_mask = buffer_1_auto_out_a_bits_mask;
	assign in_xbar_auto_in_0_a_bits_data = buffer_1_auto_out_a_bits_data;
	assign in_xbar_auto_in_0_a_bits_corrupt = buffer_1_auto_out_a_bits_corrupt;
	assign in_xbar_auto_in_0_d_ready = buffer_1_auto_out_d_ready;
	assign in_xbar_auto_out_a_ready = atomics_auto_in_a_ready;
	assign in_xbar_auto_out_d_valid = atomics_auto_in_d_valid;
	assign in_xbar_auto_out_d_bits_opcode = atomics_auto_in_d_bits_opcode;
	assign in_xbar_auto_out_d_bits_param = atomics_auto_in_d_bits_param;
	assign in_xbar_auto_out_d_bits_size = atomics_auto_in_d_bits_size;
	assign in_xbar_auto_out_d_bits_source = atomics_auto_in_d_bits_source;
	assign in_xbar_auto_out_d_bits_sink = atomics_auto_in_d_bits_sink;
	assign in_xbar_auto_out_d_bits_denied = atomics_auto_in_d_bits_denied;
	assign in_xbar_auto_out_d_bits_data = atomics_auto_in_d_bits_data;
	assign in_xbar_auto_out_d_bits_corrupt = atomics_auto_in_d_bits_corrupt;
	assign out_xbar_clock = fixedClockNode_auto_out_0_clock;
	assign out_xbar_reset = fixedClockNode_auto_out_0_reset;
	assign out_xbar_auto_in_a_valid = fixer_auto_out_a_valid;
	assign out_xbar_auto_in_a_bits_opcode = fixer_auto_out_a_bits_opcode;
	assign out_xbar_auto_in_a_bits_param = fixer_auto_out_a_bits_param;
	assign out_xbar_auto_in_a_bits_size = fixer_auto_out_a_bits_size;
	assign out_xbar_auto_in_a_bits_source = fixer_auto_out_a_bits_source;
	assign out_xbar_auto_in_a_bits_address = fixer_auto_out_a_bits_address;
	assign out_xbar_auto_in_a_bits_mask = fixer_auto_out_a_bits_mask;
	assign out_xbar_auto_in_a_bits_data = fixer_auto_out_a_bits_data;
	assign out_xbar_auto_in_a_bits_corrupt = fixer_auto_out_a_bits_corrupt;
	assign out_xbar_auto_in_d_ready = fixer_auto_out_d_ready;
	assign out_xbar_auto_out_8_a_ready = coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_ready;
	assign out_xbar_auto_out_8_d_valid = coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_valid;
	assign out_xbar_auto_out_8_d_bits_opcode = coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_opcode;
	assign out_xbar_auto_out_8_d_bits_param = coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_param;
	assign out_xbar_auto_out_8_d_bits_size = coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_size;
	assign out_xbar_auto_out_8_d_bits_source = coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_source;
	assign out_xbar_auto_out_8_d_bits_sink = coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_sink;
	assign out_xbar_auto_out_8_d_bits_denied = coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_denied;
	assign out_xbar_auto_out_8_d_bits_data = coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_data;
	assign out_xbar_auto_out_8_d_bits_corrupt = coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_bits_corrupt;
	assign out_xbar_auto_out_7_a_ready = coupler_to_slave_named_clockgater_auto_buffer_in_a_ready;
	assign out_xbar_auto_out_7_d_valid = coupler_to_slave_named_clockgater_auto_buffer_in_d_valid;
	assign out_xbar_auto_out_7_d_bits_opcode = coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_opcode;
	assign out_xbar_auto_out_7_d_bits_param = coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_param;
	assign out_xbar_auto_out_7_d_bits_size = coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_size;
	assign out_xbar_auto_out_7_d_bits_source = coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_source;
	assign out_xbar_auto_out_7_d_bits_sink = coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_sink;
	assign out_xbar_auto_out_7_d_bits_denied = coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_denied;
	assign out_xbar_auto_out_7_d_bits_data = coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_data;
	assign out_xbar_auto_out_7_d_bits_corrupt = coupler_to_slave_named_clockgater_auto_buffer_in_d_bits_corrupt;
	assign out_xbar_auto_out_6_a_ready = coupler_to_bootrom_auto_tl_in_a_ready;
	assign out_xbar_auto_out_6_d_valid = coupler_to_bootrom_auto_tl_in_d_valid;
	assign out_xbar_auto_out_6_d_bits_size = coupler_to_bootrom_auto_tl_in_d_bits_size;
	assign out_xbar_auto_out_6_d_bits_source = coupler_to_bootrom_auto_tl_in_d_bits_source;
	assign out_xbar_auto_out_6_d_bits_data = coupler_to_bootrom_auto_tl_in_d_bits_data;
	assign out_xbar_auto_out_5_a_ready = coupler_to_tile_auto_tl_in_a_ready;
	assign out_xbar_auto_out_5_d_valid = coupler_to_tile_auto_tl_in_d_valid;
	assign out_xbar_auto_out_5_d_bits_opcode = coupler_to_tile_auto_tl_in_d_bits_opcode;
	assign out_xbar_auto_out_5_d_bits_param = coupler_to_tile_auto_tl_in_d_bits_param;
	assign out_xbar_auto_out_5_d_bits_size = coupler_to_tile_auto_tl_in_d_bits_size;
	assign out_xbar_auto_out_5_d_bits_source = coupler_to_tile_auto_tl_in_d_bits_source;
	assign out_xbar_auto_out_5_d_bits_sink = coupler_to_tile_auto_tl_in_d_bits_sink;
	assign out_xbar_auto_out_5_d_bits_denied = coupler_to_tile_auto_tl_in_d_bits_denied;
	assign out_xbar_auto_out_5_d_bits_data = coupler_to_tile_auto_tl_in_d_bits_data;
	assign out_xbar_auto_out_5_d_bits_corrupt = coupler_to_tile_auto_tl_in_d_bits_corrupt;
	assign out_xbar_auto_out_4_a_ready = coupler_to_debug_auto_tl_in_a_ready;
	assign out_xbar_auto_out_4_d_valid = coupler_to_debug_auto_tl_in_d_valid;
	assign out_xbar_auto_out_4_d_bits_opcode = coupler_to_debug_auto_tl_in_d_bits_opcode;
	assign out_xbar_auto_out_4_d_bits_size = coupler_to_debug_auto_tl_in_d_bits_size;
	assign out_xbar_auto_out_4_d_bits_source = coupler_to_debug_auto_tl_in_d_bits_source;
	assign out_xbar_auto_out_4_d_bits_data = coupler_to_debug_auto_tl_in_d_bits_data;
	assign out_xbar_auto_out_3_a_ready = coupler_to_clint_auto_tl_in_a_ready;
	assign out_xbar_auto_out_3_d_valid = coupler_to_clint_auto_tl_in_d_valid;
	assign out_xbar_auto_out_3_d_bits_opcode = coupler_to_clint_auto_tl_in_d_bits_opcode;
	assign out_xbar_auto_out_3_d_bits_size = coupler_to_clint_auto_tl_in_d_bits_size;
	assign out_xbar_auto_out_3_d_bits_source = coupler_to_clint_auto_tl_in_d_bits_source;
	assign out_xbar_auto_out_3_d_bits_data = coupler_to_clint_auto_tl_in_d_bits_data;
	assign out_xbar_auto_out_2_a_ready = coupler_to_plic_auto_tl_in_a_ready;
	assign out_xbar_auto_out_2_d_valid = coupler_to_plic_auto_tl_in_d_valid;
	assign out_xbar_auto_out_2_d_bits_opcode = coupler_to_plic_auto_tl_in_d_bits_opcode;
	assign out_xbar_auto_out_2_d_bits_size = coupler_to_plic_auto_tl_in_d_bits_size;
	assign out_xbar_auto_out_2_d_bits_source = coupler_to_plic_auto_tl_in_d_bits_source;
	assign out_xbar_auto_out_2_d_bits_data = coupler_to_plic_auto_tl_in_d_bits_data;
	assign out_xbar_auto_out_1_a_ready = coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_ready;
	assign out_xbar_auto_out_1_d_valid = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_valid;
	assign out_xbar_auto_out_1_d_bits_opcode = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_opcode;
	assign out_xbar_auto_out_1_d_bits_param = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_param;
	assign out_xbar_auto_out_1_d_bits_size = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_size;
	assign out_xbar_auto_out_1_d_bits_source = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_source;
	assign out_xbar_auto_out_1_d_bits_sink = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_sink;
	assign out_xbar_auto_out_1_d_bits_denied = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_denied;
	assign out_xbar_auto_out_1_d_bits_data = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_data;
	assign out_xbar_auto_out_1_d_bits_corrupt = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_corrupt;
	assign out_xbar_auto_out_0_a_ready = wrapped_error_device_auto_buffer_in_a_ready;
	assign out_xbar_auto_out_0_d_valid = wrapped_error_device_auto_buffer_in_d_valid;
	assign out_xbar_auto_out_0_d_bits_opcode = wrapped_error_device_auto_buffer_in_d_bits_opcode;
	assign out_xbar_auto_out_0_d_bits_param = wrapped_error_device_auto_buffer_in_d_bits_param;
	assign out_xbar_auto_out_0_d_bits_size = wrapped_error_device_auto_buffer_in_d_bits_size;
	assign out_xbar_auto_out_0_d_bits_source = wrapped_error_device_auto_buffer_in_d_bits_source;
	assign out_xbar_auto_out_0_d_bits_sink = wrapped_error_device_auto_buffer_in_d_bits_sink;
	assign out_xbar_auto_out_0_d_bits_denied = wrapped_error_device_auto_buffer_in_d_bits_denied;
	assign out_xbar_auto_out_0_d_bits_data = wrapped_error_device_auto_buffer_in_d_bits_data;
	assign out_xbar_auto_out_0_d_bits_corrupt = wrapped_error_device_auto_buffer_in_d_bits_corrupt;
	assign buffer_clock = fixedClockNode_auto_out_0_clock;
	assign buffer_reset = fixedClockNode_auto_out_0_reset;
	assign buffer_auto_in_a_valid = atomics_auto_out_a_valid;
	assign buffer_auto_in_a_bits_opcode = atomics_auto_out_a_bits_opcode;
	assign buffer_auto_in_a_bits_param = atomics_auto_out_a_bits_param;
	assign buffer_auto_in_a_bits_size = atomics_auto_out_a_bits_size;
	assign buffer_auto_in_a_bits_source = atomics_auto_out_a_bits_source;
	assign buffer_auto_in_a_bits_address = atomics_auto_out_a_bits_address;
	assign buffer_auto_in_a_bits_mask = atomics_auto_out_a_bits_mask;
	assign buffer_auto_in_a_bits_data = atomics_auto_out_a_bits_data;
	assign buffer_auto_in_a_bits_corrupt = atomics_auto_out_a_bits_corrupt;
	assign buffer_auto_in_d_ready = atomics_auto_out_d_ready;
	assign buffer_auto_out_a_ready = fixer_auto_in_a_ready;
	assign buffer_auto_out_d_valid = fixer_auto_in_d_valid;
	assign buffer_auto_out_d_bits_opcode = fixer_auto_in_d_bits_opcode;
	assign buffer_auto_out_d_bits_param = fixer_auto_in_d_bits_param;
	assign buffer_auto_out_d_bits_size = fixer_auto_in_d_bits_size;
	assign buffer_auto_out_d_bits_source = fixer_auto_in_d_bits_source;
	assign buffer_auto_out_d_bits_sink = fixer_auto_in_d_bits_sink;
	assign buffer_auto_out_d_bits_denied = fixer_auto_in_d_bits_denied;
	assign buffer_auto_out_d_bits_data = fixer_auto_in_d_bits_data;
	assign buffer_auto_out_d_bits_corrupt = fixer_auto_in_d_bits_corrupt;
	assign atomics_clock = fixedClockNode_auto_out_0_clock;
	assign atomics_reset = fixedClockNode_auto_out_0_reset;
	assign atomics_auto_in_a_valid = in_xbar_auto_out_a_valid;
	assign atomics_auto_in_a_bits_opcode = in_xbar_auto_out_a_bits_opcode;
	assign atomics_auto_in_a_bits_param = in_xbar_auto_out_a_bits_param;
	assign atomics_auto_in_a_bits_size = in_xbar_auto_out_a_bits_size;
	assign atomics_auto_in_a_bits_source = in_xbar_auto_out_a_bits_source;
	assign atomics_auto_in_a_bits_address = in_xbar_auto_out_a_bits_address;
	assign atomics_auto_in_a_bits_mask = in_xbar_auto_out_a_bits_mask;
	assign atomics_auto_in_a_bits_data = in_xbar_auto_out_a_bits_data;
	assign atomics_auto_in_a_bits_corrupt = in_xbar_auto_out_a_bits_corrupt;
	assign atomics_auto_in_d_ready = in_xbar_auto_out_d_ready;
	assign atomics_auto_out_a_ready = buffer_auto_in_a_ready;
	assign atomics_auto_out_d_valid = buffer_auto_in_d_valid;
	assign atomics_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode;
	assign atomics_auto_out_d_bits_param = buffer_auto_in_d_bits_param;
	assign atomics_auto_out_d_bits_size = buffer_auto_in_d_bits_size;
	assign atomics_auto_out_d_bits_source = buffer_auto_in_d_bits_source;
	assign atomics_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink;
	assign atomics_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied;
	assign atomics_auto_out_d_bits_data = buffer_auto_in_d_bits_data;
	assign atomics_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt;
	assign wrapped_error_device_clock = fixedClockNode_auto_out_0_clock;
	assign wrapped_error_device_reset = fixedClockNode_auto_out_0_reset;
	assign wrapped_error_device_auto_buffer_in_a_valid = out_xbar_auto_out_0_a_valid;
	assign wrapped_error_device_auto_buffer_in_a_bits_opcode = out_xbar_auto_out_0_a_bits_opcode;
	assign wrapped_error_device_auto_buffer_in_a_bits_param = out_xbar_auto_out_0_a_bits_param;
	assign wrapped_error_device_auto_buffer_in_a_bits_size = out_xbar_auto_out_0_a_bits_size;
	assign wrapped_error_device_auto_buffer_in_a_bits_source = out_xbar_auto_out_0_a_bits_source;
	assign wrapped_error_device_auto_buffer_in_a_bits_address = out_xbar_auto_out_0_a_bits_address;
	assign wrapped_error_device_auto_buffer_in_a_bits_mask = out_xbar_auto_out_0_a_bits_mask;
	assign wrapped_error_device_auto_buffer_in_a_bits_corrupt = out_xbar_auto_out_0_a_bits_corrupt;
	assign wrapped_error_device_auto_buffer_in_d_ready = out_xbar_auto_out_0_d_ready;
	assign buffer_1_auto_in_a_valid = auto_bus_xing_in_a_valid;
	assign buffer_1_auto_in_a_bits_opcode = auto_bus_xing_in_a_bits_opcode;
	assign buffer_1_auto_in_a_bits_param = auto_bus_xing_in_a_bits_param;
	assign buffer_1_auto_in_a_bits_size = auto_bus_xing_in_a_bits_size;
	assign buffer_1_auto_in_a_bits_source = auto_bus_xing_in_a_bits_source;
	assign buffer_1_auto_in_a_bits_address = auto_bus_xing_in_a_bits_address;
	assign buffer_1_auto_in_a_bits_mask = auto_bus_xing_in_a_bits_mask;
	assign buffer_1_auto_in_a_bits_data = auto_bus_xing_in_a_bits_data;
	assign buffer_1_auto_in_a_bits_corrupt = auto_bus_xing_in_a_bits_corrupt;
	assign buffer_1_auto_in_d_ready = auto_bus_xing_in_d_ready;
	assign buffer_1_auto_out_a_ready = in_xbar_auto_in_0_a_ready;
	assign buffer_1_auto_out_d_valid = in_xbar_auto_in_0_d_valid;
	assign buffer_1_auto_out_d_bits_opcode = in_xbar_auto_in_0_d_bits_opcode;
	assign buffer_1_auto_out_d_bits_param = in_xbar_auto_in_0_d_bits_param;
	assign buffer_1_auto_out_d_bits_size = in_xbar_auto_in_0_d_bits_size;
	assign buffer_1_auto_out_d_bits_source = in_xbar_auto_in_0_d_bits_source;
	assign buffer_1_auto_out_d_bits_sink = in_xbar_auto_in_0_d_bits_sink;
	assign buffer_1_auto_out_d_bits_denied = in_xbar_auto_in_0_d_bits_denied;
	assign buffer_1_auto_out_d_bits_data = in_xbar_auto_in_0_d_bits_data;
	assign buffer_1_auto_out_d_bits_corrupt = in_xbar_auto_in_0_d_bits_corrupt;
	assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_valid = out_xbar_auto_out_1_a_valid;
	assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_opcode = out_xbar_auto_out_1_a_bits_opcode;
	assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_param = out_xbar_auto_out_1_a_bits_param;
	assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_size = out_xbar_auto_out_1_a_bits_size;
	assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_source = out_xbar_auto_out_1_a_bits_source;
	assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_address = out_xbar_auto_out_1_a_bits_address;
	assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_mask = out_xbar_auto_out_1_a_bits_mask;
	assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_data = out_xbar_auto_out_1_a_bits_data;
	assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_corrupt = out_xbar_auto_out_1_a_bits_corrupt;
	assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_ready = out_xbar_auto_out_1_d_ready;
	assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_ready = auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready;
	assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_valid = auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid;
	assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_opcode = auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode;
	assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_param = auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_param;
	assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_size = auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size;
	assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_source = auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source;
	assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_sink = auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_sink;
	assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_denied = auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied;
	assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_data = auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data;
	assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_corrupt = auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt;
	assign coupler_to_plic_clock = fixedClockNode_auto_out_0_clock;
	assign coupler_to_plic_reset = fixedClockNode_auto_out_0_reset;
	assign coupler_to_plic_auto_fragmenter_out_a_ready = auto_coupler_to_plic_fragmenter_out_a_ready;
	assign coupler_to_plic_auto_fragmenter_out_d_valid = auto_coupler_to_plic_fragmenter_out_d_valid;
	assign coupler_to_plic_auto_fragmenter_out_d_bits_opcode = auto_coupler_to_plic_fragmenter_out_d_bits_opcode;
	assign coupler_to_plic_auto_fragmenter_out_d_bits_size = auto_coupler_to_plic_fragmenter_out_d_bits_size;
	assign coupler_to_plic_auto_fragmenter_out_d_bits_source = auto_coupler_to_plic_fragmenter_out_d_bits_source;
	assign coupler_to_plic_auto_fragmenter_out_d_bits_data = auto_coupler_to_plic_fragmenter_out_d_bits_data;
	assign coupler_to_plic_auto_tl_in_a_valid = out_xbar_auto_out_2_a_valid;
	assign coupler_to_plic_auto_tl_in_a_bits_opcode = out_xbar_auto_out_2_a_bits_opcode;
	assign coupler_to_plic_auto_tl_in_a_bits_param = out_xbar_auto_out_2_a_bits_param;
	assign coupler_to_plic_auto_tl_in_a_bits_size = out_xbar_auto_out_2_a_bits_size;
	assign coupler_to_plic_auto_tl_in_a_bits_source = out_xbar_auto_out_2_a_bits_source;
	assign coupler_to_plic_auto_tl_in_a_bits_address = out_xbar_auto_out_2_a_bits_address;
	assign coupler_to_plic_auto_tl_in_a_bits_mask = out_xbar_auto_out_2_a_bits_mask;
	assign coupler_to_plic_auto_tl_in_a_bits_data = out_xbar_auto_out_2_a_bits_data;
	assign coupler_to_plic_auto_tl_in_a_bits_corrupt = out_xbar_auto_out_2_a_bits_corrupt;
	assign coupler_to_plic_auto_tl_in_d_ready = out_xbar_auto_out_2_d_ready;
	assign coupler_to_clint_clock = fixedClockNode_auto_out_0_clock;
	assign coupler_to_clint_reset = fixedClockNode_auto_out_0_reset;
	assign coupler_to_clint_auto_fragmenter_out_a_ready = auto_coupler_to_clint_fragmenter_out_a_ready;
	assign coupler_to_clint_auto_fragmenter_out_d_valid = auto_coupler_to_clint_fragmenter_out_d_valid;
	assign coupler_to_clint_auto_fragmenter_out_d_bits_opcode = auto_coupler_to_clint_fragmenter_out_d_bits_opcode;
	assign coupler_to_clint_auto_fragmenter_out_d_bits_size = auto_coupler_to_clint_fragmenter_out_d_bits_size;
	assign coupler_to_clint_auto_fragmenter_out_d_bits_source = auto_coupler_to_clint_fragmenter_out_d_bits_source;
	assign coupler_to_clint_auto_fragmenter_out_d_bits_data = auto_coupler_to_clint_fragmenter_out_d_bits_data;
	assign coupler_to_clint_auto_tl_in_a_valid = out_xbar_auto_out_3_a_valid;
	assign coupler_to_clint_auto_tl_in_a_bits_opcode = out_xbar_auto_out_3_a_bits_opcode;
	assign coupler_to_clint_auto_tl_in_a_bits_param = out_xbar_auto_out_3_a_bits_param;
	assign coupler_to_clint_auto_tl_in_a_bits_size = out_xbar_auto_out_3_a_bits_size;
	assign coupler_to_clint_auto_tl_in_a_bits_source = out_xbar_auto_out_3_a_bits_source;
	assign coupler_to_clint_auto_tl_in_a_bits_address = out_xbar_auto_out_3_a_bits_address;
	assign coupler_to_clint_auto_tl_in_a_bits_mask = out_xbar_auto_out_3_a_bits_mask;
	assign coupler_to_clint_auto_tl_in_a_bits_data = out_xbar_auto_out_3_a_bits_data;
	assign coupler_to_clint_auto_tl_in_a_bits_corrupt = out_xbar_auto_out_3_a_bits_corrupt;
	assign coupler_to_clint_auto_tl_in_d_ready = out_xbar_auto_out_3_d_ready;
	assign coupler_to_debug_clock = fixedClockNode_auto_out_0_clock;
	assign coupler_to_debug_reset = fixedClockNode_auto_out_0_reset;
	assign coupler_to_debug_auto_fragmenter_out_a_ready = auto_coupler_to_debug_fragmenter_out_a_ready;
	assign coupler_to_debug_auto_fragmenter_out_d_valid = auto_coupler_to_debug_fragmenter_out_d_valid;
	assign coupler_to_debug_auto_fragmenter_out_d_bits_opcode = auto_coupler_to_debug_fragmenter_out_d_bits_opcode;
	assign coupler_to_debug_auto_fragmenter_out_d_bits_size = auto_coupler_to_debug_fragmenter_out_d_bits_size;
	assign coupler_to_debug_auto_fragmenter_out_d_bits_source = auto_coupler_to_debug_fragmenter_out_d_bits_source;
	assign coupler_to_debug_auto_fragmenter_out_d_bits_data = auto_coupler_to_debug_fragmenter_out_d_bits_data;
	assign coupler_to_debug_auto_tl_in_a_valid = out_xbar_auto_out_4_a_valid;
	assign coupler_to_debug_auto_tl_in_a_bits_opcode = out_xbar_auto_out_4_a_bits_opcode;
	assign coupler_to_debug_auto_tl_in_a_bits_param = out_xbar_auto_out_4_a_bits_param;
	assign coupler_to_debug_auto_tl_in_a_bits_size = out_xbar_auto_out_4_a_bits_size;
	assign coupler_to_debug_auto_tl_in_a_bits_source = out_xbar_auto_out_4_a_bits_source;
	assign coupler_to_debug_auto_tl_in_a_bits_address = out_xbar_auto_out_4_a_bits_address;
	assign coupler_to_debug_auto_tl_in_a_bits_mask = out_xbar_auto_out_4_a_bits_mask;
	assign coupler_to_debug_auto_tl_in_a_bits_data = out_xbar_auto_out_4_a_bits_data;
	assign coupler_to_debug_auto_tl_in_a_bits_corrupt = out_xbar_auto_out_4_a_bits_corrupt;
	assign coupler_to_debug_auto_tl_in_d_ready = out_xbar_auto_out_4_d_ready;
	assign coupler_to_tile_auto_tl_slave_clock_xing_out_a_ready = auto_coupler_to_tile_tl_slave_clock_xing_out_a_ready;
	assign coupler_to_tile_auto_tl_slave_clock_xing_out_d_valid = auto_coupler_to_tile_tl_slave_clock_xing_out_d_valid;
	assign coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_opcode = auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_opcode;
	assign coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_param = auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_param;
	assign coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_size = auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_size;
	assign coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_source = auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_source;
	assign coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_sink = auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_sink;
	assign coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_denied = auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_denied;
	assign coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_data = auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_data;
	assign coupler_to_tile_auto_tl_slave_clock_xing_out_d_bits_corrupt = auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_corrupt;
	assign coupler_to_tile_auto_tl_in_a_valid = out_xbar_auto_out_5_a_valid;
	assign coupler_to_tile_auto_tl_in_a_bits_opcode = out_xbar_auto_out_5_a_bits_opcode;
	assign coupler_to_tile_auto_tl_in_a_bits_param = out_xbar_auto_out_5_a_bits_param;
	assign coupler_to_tile_auto_tl_in_a_bits_size = out_xbar_auto_out_5_a_bits_size;
	assign coupler_to_tile_auto_tl_in_a_bits_source = out_xbar_auto_out_5_a_bits_source;
	assign coupler_to_tile_auto_tl_in_a_bits_address = out_xbar_auto_out_5_a_bits_address;
	assign coupler_to_tile_auto_tl_in_a_bits_mask = out_xbar_auto_out_5_a_bits_mask;
	assign coupler_to_tile_auto_tl_in_a_bits_data = out_xbar_auto_out_5_a_bits_data;
	assign coupler_to_tile_auto_tl_in_d_ready = out_xbar_auto_out_5_d_ready;
	assign coupler_to_bootrom_clock = fixedClockNode_auto_out_0_clock;
	assign coupler_to_bootrom_reset = fixedClockNode_auto_out_0_reset;
	assign coupler_to_bootrom_auto_fragmenter_out_a_ready = auto_coupler_to_bootrom_fragmenter_out_a_ready;
	assign coupler_to_bootrom_auto_fragmenter_out_d_valid = auto_coupler_to_bootrom_fragmenter_out_d_valid;
	assign coupler_to_bootrom_auto_fragmenter_out_d_bits_size = auto_coupler_to_bootrom_fragmenter_out_d_bits_size;
	assign coupler_to_bootrom_auto_fragmenter_out_d_bits_source = auto_coupler_to_bootrom_fragmenter_out_d_bits_source;
	assign coupler_to_bootrom_auto_fragmenter_out_d_bits_data = auto_coupler_to_bootrom_fragmenter_out_d_bits_data;
	assign coupler_to_bootrom_auto_tl_in_a_valid = out_xbar_auto_out_6_a_valid;
	assign coupler_to_bootrom_auto_tl_in_a_bits_opcode = out_xbar_auto_out_6_a_bits_opcode;
	assign coupler_to_bootrom_auto_tl_in_a_bits_param = out_xbar_auto_out_6_a_bits_param;
	assign coupler_to_bootrom_auto_tl_in_a_bits_size = out_xbar_auto_out_6_a_bits_size;
	assign coupler_to_bootrom_auto_tl_in_a_bits_source = out_xbar_auto_out_6_a_bits_source;
	assign coupler_to_bootrom_auto_tl_in_a_bits_address = out_xbar_auto_out_6_a_bits_address;
	assign coupler_to_bootrom_auto_tl_in_a_bits_mask = out_xbar_auto_out_6_a_bits_mask;
	assign coupler_to_bootrom_auto_tl_in_a_bits_corrupt = out_xbar_auto_out_6_a_bits_corrupt;
	assign coupler_to_bootrom_auto_tl_in_d_ready = out_xbar_auto_out_6_d_ready;
	assign coupler_from_port_named_custom_boot_pin_auto_tl_in_a_valid = (3'h0 == state ? 1'h0 : _GEN_28);
	assign coupler_from_port_named_custom_boot_pin_auto_tl_in_a_bits_address = (3'h1 == state ? 32'h00004000 : 32'h02000000);
	assign coupler_from_port_named_custom_boot_pin_auto_tl_in_a_bits_data = (3'h1 == state ? 32'h80000000 : 32'h00000001);
	assign coupler_from_port_named_custom_boot_pin_auto_tl_out_a_ready = in_xbar_auto_in_1_a_ready;
	assign coupler_from_port_named_custom_boot_pin_auto_tl_out_d_valid = in_xbar_auto_in_1_d_valid;
	assign coupler_to_slave_named_clockgater_clock = fixedClockNode_auto_out_0_clock;
	assign coupler_to_slave_named_clockgater_reset = fixedClockNode_auto_out_0_reset;
	assign coupler_to_slave_named_clockgater_auto_buffer_in_a_valid = out_xbar_auto_out_7_a_valid;
	assign coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_opcode = out_xbar_auto_out_7_a_bits_opcode;
	assign coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_param = out_xbar_auto_out_7_a_bits_param;
	assign coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_size = out_xbar_auto_out_7_a_bits_size;
	assign coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_source = out_xbar_auto_out_7_a_bits_source;
	assign coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_address = out_xbar_auto_out_7_a_bits_address;
	assign coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_mask = out_xbar_auto_out_7_a_bits_mask;
	assign coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_data = out_xbar_auto_out_7_a_bits_data;
	assign coupler_to_slave_named_clockgater_auto_buffer_in_a_bits_corrupt = out_xbar_auto_out_7_a_bits_corrupt;
	assign coupler_to_slave_named_clockgater_auto_buffer_in_d_ready = out_xbar_auto_out_7_d_ready;
	assign coupler_to_slave_named_clockgater_auto_buffer_out_a_ready = auto_coupler_to_slave_named_clockgater_buffer_out_a_ready;
	assign coupler_to_slave_named_clockgater_auto_buffer_out_d_valid = auto_coupler_to_slave_named_clockgater_buffer_out_d_valid;
	assign coupler_to_slave_named_clockgater_auto_buffer_out_d_bits_opcode = auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_opcode;
	assign coupler_to_slave_named_clockgater_auto_buffer_out_d_bits_size = auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_size;
	assign coupler_to_slave_named_clockgater_auto_buffer_out_d_bits_source = auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_source;
	assign coupler_to_slave_named_clockgater_auto_buffer_out_d_bits_data = auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_data;
	assign coupler_to_slave_named_tileresetsetter_clock = fixedClockNode_auto_out_0_clock;
	assign coupler_to_slave_named_tileresetsetter_reset = fixedClockNode_auto_out_0_reset;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_valid = out_xbar_auto_out_8_a_valid;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_opcode = out_xbar_auto_out_8_a_bits_opcode;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_param = out_xbar_auto_out_8_a_bits_param;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_size = out_xbar_auto_out_8_a_bits_size;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_source = out_xbar_auto_out_8_a_bits_source;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_address = out_xbar_auto_out_8_a_bits_address;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_mask = out_xbar_auto_out_8_a_bits_mask;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_data = out_xbar_auto_out_8_a_bits_data;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_in_a_bits_corrupt = out_xbar_auto_out_8_a_bits_corrupt;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_in_d_ready = out_xbar_auto_out_8_d_ready;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_out_a_ready = auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_ready;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_valid = auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_valid;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_bits_opcode = auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_opcode;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_bits_size = auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_size;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_bits_source = auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_source;
	assign coupler_to_slave_named_tileresetsetter_auto_buffer_out_d_bits_data = auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_data;
	always @(posedge bundleIn_0_clock)
		if (bundleIn_0_reset)
			state <= 3'h0;
		else if (3'h0 == state) begin
			if (custom_boot)
				state <= 3'h1;
		end
		else if (3'h1 == state) begin
			if (_T_2)
				state <= 3'h2;
		end
		else if (3'h2 == state)
			state <= _GEN_2;
		else
			state <= _GEN_17;
endmodule
module TLMonitor_31 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_15 = io_in_a_bits_opcode == 3'h6;
	wire _T_17 = io_in_a_bits_size <= 4'hc;
	wire [32:0] _T_26 = $signed(_T_7) & -33'sh000005000;
	wire _T_27 = $signed(_T_26) == 33'sh000000000;
	wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_29 = {1'b0, $signed(_T_28)};
	wire [32:0] _T_31 = $signed(_T_29) & -33'sh000001000;
	wire _T_32 = $signed(_T_31) == 33'sh000000000;
	wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [32:0] _T_36 = $signed(_T_34) & -33'sh000010000;
	wire _T_37 = $signed(_T_36) == 33'sh000000000;
	wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_39 = {1'b0, $signed(_T_38)};
	wire [32:0] _T_41 = $signed(_T_39) & -33'sh000010000;
	wire _T_42 = $signed(_T_41) == 33'sh000000000;
	wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_44 = {1'b0, $signed(_T_43)};
	wire [32:0] _T_46 = $signed(_T_44) & -33'sh000011000;
	wire _T_47 = $signed(_T_46) == 33'sh000000000;
	wire [31:0] _T_48 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_49 = {1'b0, $signed(_T_48)};
	wire [32:0] _T_51 = $signed(_T_49) & -33'sh000010000;
	wire _T_52 = $signed(_T_51) == 33'sh000000000;
	wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_54 = {1'b0, $signed(_T_53)};
	wire [32:0] _T_56 = $signed(_T_54) & -33'sh004000000;
	wire _T_57 = $signed(_T_56) == 33'sh000000000;
	wire [31:0] _T_58 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_59 = {1'b0, $signed(_T_58)};
	wire [32:0] _T_61 = $signed(_T_59) & -33'sh000001000;
	wire _T_62 = $signed(_T_61) == 33'sh000000000;
	wire [31:0] _T_63 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_64 = {1'b0, $signed(_T_63)};
	wire [32:0] _T_66 = $signed(_T_64) & -33'sh000001000;
	wire _T_67 = $signed(_T_66) == 33'sh000000000;
	wire [31:0] _T_68 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_69 = {1'b0, $signed(_T_68)};
	wire [32:0] _T_71 = $signed(_T_69) & -33'sh000004000;
	wire _T_72 = $signed(_T_71) == 33'sh000000000;
	wire _T_167 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_171 = ~io_in_a_bits_mask;
	wire _T_172 = _T_171 == 4'h0;
	wire _T_180 = io_in_a_bits_opcode == 3'h7;
	wire _T_336 = io_in_a_bits_param != 3'h0;
	wire _T_349 = io_in_a_bits_opcode == 3'h4;
	wire _T_368 = _T_17 & _T_32;
	wire _T_370 = io_in_a_bits_size <= 4'h6;
	wire _T_425 = (((((((_T_27 | _T_37) | _T_42) | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_426 = _T_370 & _T_425;
	wire _T_428 = _T_368 | _T_426;
	wire _T_438 = io_in_a_bits_param == 3'h0;
	wire _T_442 = io_in_a_bits_mask == mask;
	wire _T_450 = io_in_a_bits_opcode == 3'h0;
	wire _T_511 = (((((_T_27 | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_512 = _T_370 & _T_511;
	wire _T_527 = _T_368 | _T_512;
	wire _T_529 = _T_17 & _T_527;
	wire _T_547 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_640 = ~mask;
	wire [3:0] _T_641 = io_in_a_bits_mask & _T_640;
	wire _T_642 = _T_641 == 4'h0;
	wire _T_646 = io_in_a_bits_opcode == 3'h2;
	wire _T_654 = io_in_a_bits_size <= 4'h2;
	wire _T_703 = ((((((_T_27 | _T_32) | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_704 = _T_654 & _T_703;
	wire _T_720 = _T_17 & _T_704;
	wire _T_730 = io_in_a_bits_param <= 3'h4;
	wire _T_738 = io_in_a_bits_opcode == 3'h3;
	wire _T_822 = io_in_a_bits_param <= 3'h3;
	wire _T_830 = io_in_a_bits_opcode == 3'h5;
	wire _T_904 = _T_17 & _T_368;
	wire _T_914 = io_in_a_bits_param <= 3'h1;
	wire _T_926 = io_in_d_bits_opcode <= 3'h6;
	wire _T_930 = io_in_d_bits_opcode == 3'h6;
	wire _T_934 = io_in_d_bits_size >= 4'h2;
	wire _T_938 = io_in_d_bits_param == 2'h0;
	wire _T_942 = ~io_in_d_bits_corrupt;
	wire _T_946 = ~io_in_d_bits_denied;
	wire _T_950 = io_in_d_bits_opcode == 3'h4;
	wire _T_961 = io_in_d_bits_param <= 2'h2;
	wire _T_965 = io_in_d_bits_param != 2'h2;
	wire _T_978 = io_in_d_bits_opcode == 3'h5;
	wire _T_998 = _T_946 | io_in_d_bits_corrupt;
	wire _T_1007 = io_in_d_bits_opcode == 3'h0;
	wire _T_1024 = io_in_d_bits_opcode == 3'h1;
	wire _T_1042 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg [31:0] address;
	wire _T_1072 = io_in_a_valid & ~a_first;
	wire _T_1073 = io_in_a_bits_opcode == opcode;
	wire _T_1077 = io_in_a_bits_param == param;
	wire _T_1081 = io_in_a_bits_size == size;
	wire _T_1089 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg sink;
	reg denied;
	wire _T_1096 = io_in_d_valid & ~d_first;
	wire _T_1097 = io_in_d_bits_opcode == opcode_1;
	wire _T_1101 = io_in_d_bits_param == param_1;
	wire _T_1105 = io_in_d_bits_size == size_1;
	wire _T_1113 = io_in_d_bits_sink == sink;
	wire _T_1117 = io_in_d_bits_denied == denied;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [7:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_72 = {12'd0, inflight_opcodes};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_72 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [15:0] _GEN_74 = {8'd0, inflight_sizes};
	wire [15:0] _a_size_lookup_T_6 = _GEN_74 & _a_size_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_1123 = io_in_a_valid & a_first_1;
	wire [1:0] _GEN_15 = (io_in_a_valid & a_first_1 ? 2'h1 : 2'h0);
	wire _T_1126 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _a_opcodes_set_T_1 = {15'd0, a_opcodes_set_interm};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [19:0] _a_sizes_set_T_1 = {15'd0, a_sizes_set_interm};
	wire _T_1130 = ~inflight;
	wire [1:0] _GEN_16 = (_a_first_T & a_first_1 ? 2'h1 : 2'h0);
	wire [18:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [19:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 20'h00000);
	wire _T_1134 = io_in_d_valid & d_first_1;
	wire _T_1136 = ~_T_930;
	wire _T_1137 = (io_in_d_valid & d_first_1) & ~_T_930;
	wire [1:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_930 ? 2'h1 : 2'h0);
	wire [30:0] _d_opcodes_clr_T_5 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_sizes_clr_T_5 = {15'd0, _a_size_lookup_T_5};
	wire [1:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_1136 ? 2'h1 : 2'h0);
	wire [30:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1136 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [30:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1136 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire _T_1149 = inflight | _T_1123;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1154 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1155 = (io_in_d_bits_opcode == _GEN_32) | _T_1154;
	wire _T_1159 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1166 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1167 = (io_in_d_bits_opcode == _GEN_48) | _T_1166;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_76 = {4'd0, io_in_d_bits_size};
	wire _T_1171 = _GEN_76 == a_size_lookup;
	wire _T_1181 = ((_T_1134 & a_first_1) & io_in_a_valid) & _T_1136;
	wire _T_1183 = ~io_in_d_ready | io_in_a_ready;
	wire a_set_wo_ready = _GEN_15[0];
	wire d_clr_wo_ready = _GEN_21[0];
	wire _T_1190 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire a_set = _GEN_16[0];
	wire d_clr = _GEN_22[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [7:0] a_sizes_set = _GEN_20[7:0];
	wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [7:0] d_sizes_clr = _GEN_24[7:0];
	wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1199 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [7:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [15:0] _GEN_79 = {8'd0, inflight_sizes_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_79 & _a_size_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_1225 = (io_in_d_valid & d_first_2) & _T_930;
	wire [30:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_930 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1243 = _GEN_76 == c_size_lookup;
	wire [7:0] d_sizes_clr_1 = _GEN_69[7:0];
	wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 8'h00;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 8'h00;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module TLMonitor_32 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_address,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [31:0] io_in_a_bits_address;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire [31:0] _is_aligned_T = io_in_a_bits_address & 32'h0000003f;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire [32:0] _T_26 = $signed(_T_7) & -33'sh000005000;
	wire _T_27 = $signed(_T_26) == 33'sh000000000;
	wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_29 = {1'b0, $signed(_T_28)};
	wire [32:0] _T_31 = $signed(_T_29) & -33'sh000001000;
	wire _T_32 = $signed(_T_31) == 33'sh000000000;
	wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [32:0] _T_36 = $signed(_T_34) & -33'sh000010000;
	wire _T_37 = $signed(_T_36) == 33'sh000000000;
	wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_39 = {1'b0, $signed(_T_38)};
	wire [32:0] _T_41 = $signed(_T_39) & -33'sh000010000;
	wire _T_42 = $signed(_T_41) == 33'sh000000000;
	wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_44 = {1'b0, $signed(_T_43)};
	wire [32:0] _T_46 = $signed(_T_44) & -33'sh000011000;
	wire _T_47 = $signed(_T_46) == 33'sh000000000;
	wire [31:0] _T_48 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_49 = {1'b0, $signed(_T_48)};
	wire [32:0] _T_51 = $signed(_T_49) & -33'sh000010000;
	wire _T_52 = $signed(_T_51) == 33'sh000000000;
	wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_54 = {1'b0, $signed(_T_53)};
	wire [32:0] _T_56 = $signed(_T_54) & -33'sh004000000;
	wire _T_57 = $signed(_T_56) == 33'sh000000000;
	wire [31:0] _T_58 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_59 = {1'b0, $signed(_T_58)};
	wire [32:0] _T_61 = $signed(_T_59) & -33'sh000001000;
	wire _T_62 = $signed(_T_61) == 33'sh000000000;
	wire [31:0] _T_63 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_64 = {1'b0, $signed(_T_63)};
	wire [32:0] _T_66 = $signed(_T_64) & -33'sh000001000;
	wire _T_67 = $signed(_T_66) == 33'sh000000000;
	wire [31:0] _T_68 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_69 = {1'b0, $signed(_T_68)};
	wire [32:0] _T_71 = $signed(_T_69) & -33'sh000004000;
	wire _T_72 = $signed(_T_71) == 33'sh000000000;
	wire _T_425 = (((((((_T_27 | _T_37) | _T_42) | _T_47) | _T_52) | _T_57) | _T_62) | _T_67) | _T_72;
	wire _T_428 = _T_32 | _T_425;
	wire _T_926 = io_in_d_bits_opcode <= 3'h6;
	wire _T_930 = io_in_d_bits_opcode == 3'h6;
	wire _T_934 = io_in_d_bits_size >= 4'h2;
	wire _T_938 = io_in_d_bits_param == 2'h0;
	wire _T_942 = ~io_in_d_bits_corrupt;
	wire _T_946 = ~io_in_d_bits_denied;
	wire _T_950 = io_in_d_bits_opcode == 3'h4;
	wire _T_961 = io_in_d_bits_param <= 2'h2;
	wire _T_965 = io_in_d_bits_param != 2'h2;
	wire _T_978 = io_in_d_bits_opcode == 3'h5;
	wire _T_998 = _T_946 | io_in_d_bits_corrupt;
	wire _T_1007 = io_in_d_bits_opcode == 3'h0;
	wire _T_1024 = io_in_d_bits_opcode == 3'h1;
	wire _T_1042 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [31:0] address;
	wire _T_1072 = io_in_a_valid & ~a_first;
	wire _T_1089 = io_in_a_bits_address == address;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg sink;
	reg denied;
	wire _T_1096 = io_in_d_valid & ~d_first;
	wire _T_1097 = io_in_d_bits_opcode == opcode_1;
	wire _T_1101 = io_in_d_bits_param == param_1;
	wire _T_1105 = io_in_d_bits_size == size_1;
	wire _T_1113 = io_in_d_bits_sink == sink;
	wire _T_1117 = io_in_d_bits_denied == denied;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [7:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_71 = {12'd0, inflight_opcodes};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_71 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [15:0] _GEN_73 = {8'd0, inflight_sizes};
	wire [15:0] _a_size_lookup_T_6 = _GEN_73 & _a_size_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_1123 = io_in_a_valid & a_first_1;
	wire [1:0] _GEN_15 = (io_in_a_valid & a_first_1 ? 2'h1 : 2'h0);
	wire _T_1126 = a_first_done & a_first_1;
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? 4'h9 : 4'h0);
	wire [18:0] _a_opcodes_set_T_1 = {15'd0, a_opcodes_set_interm};
	wire [4:0] a_sizes_set_interm = (a_first_done & a_first_1 ? 5'h0d : 5'h00);
	wire [19:0] _a_sizes_set_T_1 = {15'd0, a_sizes_set_interm};
	wire _T_1130 = ~inflight;
	wire [1:0] _GEN_16 = (a_first_done & a_first_1 ? 2'h1 : 2'h0);
	wire [18:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [19:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 20'h00000);
	wire _T_1134 = io_in_d_valid & d_first_1;
	wire _T_1136 = ~_T_930;
	wire _T_1137 = (io_in_d_valid & d_first_1) & ~_T_930;
	wire [1:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_930 ? 2'h1 : 2'h0);
	wire [30:0] _d_opcodes_clr_T_5 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_sizes_clr_T_5 = {15'd0, _a_size_lookup_T_5};
	wire [30:0] _GEN_23 = (_T_1137 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [30:0] _GEN_24 = (_T_1137 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire _T_1149 = inflight | _T_1123;
	wire _T_1155 = _T_1024 | _T_1024;
	wire _T_1159 = 4'h6 == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1166 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1167 = (io_in_d_bits_opcode == _GEN_48) | _T_1166;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_75 = {4'd0, io_in_d_bits_size};
	wire _T_1171 = _GEN_75 == a_size_lookup;
	wire _T_1181 = ((_T_1134 & a_first_1) & io_in_a_valid) & _T_1136;
	wire a_set_wo_ready = _GEN_15[0];
	wire d_clr_wo_ready = _GEN_21[0];
	wire _T_1190 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire a_set = _GEN_16[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [7:0] a_sizes_set = _GEN_20[7:0];
	wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [7:0] d_sizes_clr = _GEN_24[7:0];
	wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1199 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [7:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [15:0] _GEN_78 = {8'd0, inflight_sizes_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_78 & _a_size_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_1225 = (io_in_d_valid & d_first_2) & _T_930;
	wire [30:0] _GEN_69 = (_T_1225 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1243 = _GEN_75 == c_size_lookup;
	wire [7:0] d_sizes_clr_1 = _GEN_69[7:0];
	wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 10'h000;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (io_in_d_valid)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (io_in_d_valid & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (io_in_d_valid & d_first)
			param_1 <= io_in_d_bits_param;
		if (io_in_d_valid & d_first)
			size_1 <= io_in_d_bits_size;
		if (io_in_d_valid & d_first)
			sink <= io_in_d_bits_sink;
		if (io_in_d_valid & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr_wo_ready;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 8'h00;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 10'h000;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (io_in_d_valid)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | io_in_d_valid)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 8'h00;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (io_in_d_valid)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module TLXbar_6 (
	clock,
	reset,
	auto_in_1_a_ready,
	auto_in_1_a_valid,
	auto_in_1_a_bits_address,
	auto_in_1_d_valid,
	auto_in_1_d_bits_opcode,
	auto_in_1_d_bits_size,
	auto_in_1_d_bits_data,
	auto_in_1_d_bits_corrupt,
	auto_in_0_a_ready,
	auto_in_0_a_valid,
	auto_in_0_a_bits_opcode,
	auto_in_0_a_bits_param,
	auto_in_0_a_bits_size,
	auto_in_0_a_bits_address,
	auto_in_0_a_bits_mask,
	auto_in_0_a_bits_data,
	auto_in_0_d_ready,
	auto_in_0_d_valid,
	auto_in_0_d_bits_opcode,
	auto_in_0_d_bits_size,
	auto_in_0_d_bits_denied,
	auto_in_0_d_bits_data,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_1_a_ready;
	input auto_in_1_a_valid;
	input [31:0] auto_in_1_a_bits_address;
	output wire auto_in_1_d_valid;
	output wire [2:0] auto_in_1_d_bits_opcode;
	output wire [3:0] auto_in_1_d_bits_size;
	output wire [31:0] auto_in_1_d_bits_data;
	output wire auto_in_1_d_bits_corrupt;
	output wire auto_in_0_a_ready;
	input auto_in_0_a_valid;
	input [2:0] auto_in_0_a_bits_opcode;
	input [2:0] auto_in_0_a_bits_param;
	input [3:0] auto_in_0_a_bits_size;
	input [31:0] auto_in_0_a_bits_address;
	input [3:0] auto_in_0_a_bits_mask;
	input [31:0] auto_in_0_a_bits_data;
	input auto_in_0_d_ready;
	output wire auto_in_0_d_valid;
	output wire [2:0] auto_in_0_d_bits_opcode;
	output wire [3:0] auto_in_0_d_bits_size;
	output wire auto_in_0_d_bits_denied;
	output wire [31:0] auto_in_0_d_bits_data;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire [31:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [3:0] monitor_io_in_d_bits_size;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire monitor_1_clock;
	wire monitor_1_reset;
	wire monitor_1_io_in_a_ready;
	wire monitor_1_io_in_a_valid;
	wire [31:0] monitor_1_io_in_a_bits_address;
	wire monitor_1_io_in_d_valid;
	wire [2:0] monitor_1_io_in_d_bits_opcode;
	wire [1:0] monitor_1_io_in_d_bits_param;
	wire [3:0] monitor_1_io_in_d_bits_size;
	wire monitor_1_io_in_d_bits_sink;
	wire monitor_1_io_in_d_bits_denied;
	wire monitor_1_io_in_d_bits_corrupt;
	wire requestDOI_0_1 = ~auto_out_d_bits_source;
	wire [26:0] _beatsAI_decode_T_1 = 27'h0000fff << auto_in_0_a_bits_size;
	wire [11:0] _beatsAI_decode_T_3 = ~_beatsAI_decode_T_1[11:0];
	wire [9:0] beatsAI_decode = _beatsAI_decode_T_3[11:2];
	wire beatsAI_opdata = ~auto_in_0_a_bits_opcode[2];
	reg [9:0] beatsLeft;
	wire idle = beatsLeft == 10'h000;
	wire latch = idle & auto_out_a_ready;
	wire [1:0] readys_valid = {auto_in_1_a_valid, auto_in_0_a_valid};
	wire _readys_T_3 = ~reset;
	reg [1:0] readys_mask;
	wire [1:0] _readys_filter_T = ~readys_mask;
	wire [1:0] _readys_filter_T_1 = readys_valid & _readys_filter_T;
	wire [3:0] readys_filter = {_readys_filter_T_1, auto_in_1_a_valid, auto_in_0_a_valid};
	wire [3:0] _GEN_1 = {1'd0, readys_filter[3:1]};
	wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_1;
	wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0};
	wire [3:0] _GEN_2 = {1'd0, _readys_unready_T_1[3:1]};
	wire [3:0] readys_unready = _GEN_2 | _readys_unready_T_4;
	wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0];
	wire [1:0] readys_readys = ~_readys_readys_T_2;
	wire [1:0] _readys_mask_T = readys_readys & readys_valid;
	wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0};
	wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0];
	wire readys_0 = readys_readys[0];
	wire readys_1 = readys_readys[1];
	wire earlyWinner_0 = readys_0 & auto_in_0_a_valid;
	wire earlyWinner_1 = readys_1 & auto_in_1_a_valid;
	wire _prefixOR_T = earlyWinner_0 | earlyWinner_1;
	wire _T_10 = auto_in_0_a_valid | auto_in_1_a_valid;
	wire _T_11 = ~(auto_in_0_a_valid | auto_in_1_a_valid);
	reg state_0;
	wire muxStateEarly_0 = (idle ? earlyWinner_0 : state_0);
	reg state_1;
	wire muxStateEarly_1 = (idle ? earlyWinner_1 : state_1);
	wire _out_0_a_earlyValid_T_3 = (state_0 & auto_in_0_a_valid) | (state_1 & auto_in_1_a_valid);
	wire out_2_0_a_earlyValid = (idle ? _T_10 : _out_0_a_earlyValid_T_3);
	wire _beatsLeft_T_2 = auto_out_a_ready & out_2_0_a_earlyValid;
	wire [9:0] _GEN_3 = {9'd0, _beatsLeft_T_2};
	wire [9:0] _beatsLeft_T_4 = beatsLeft - _GEN_3;
	wire allowed_0 = (idle ? readys_0 : state_0);
	wire allowed_1 = (idle ? readys_1 : state_1);
	wire [3:0] _T_30 = (muxStateEarly_0 ? auto_in_0_a_bits_mask : 4'h0);
	wire [3:0] _T_31 = (muxStateEarly_1 ? 4'hf : 4'h0);
	wire [31:0] _T_33 = (muxStateEarly_0 ? auto_in_0_a_bits_address : 32'h00000000);
	wire [31:0] _T_34 = (muxStateEarly_1 ? auto_in_1_a_bits_address : 32'h00000000);
	wire [3:0] _T_39 = (muxStateEarly_0 ? auto_in_0_a_bits_size : 4'h0);
	wire [3:0] _T_40 = (muxStateEarly_1 ? 4'h6 : 4'h0);
	wire [2:0] _T_45 = (muxStateEarly_0 ? auto_in_0_a_bits_opcode : 3'h0);
	wire [2:0] _T_46 = (muxStateEarly_1 ? 3'h4 : 3'h0);
	TLMonitor_31 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	TLMonitor_32 monitor_1(
		.clock(monitor_1_clock),
		.reset(monitor_1_reset),
		.io_in_a_ready(monitor_1_io_in_a_ready),
		.io_in_a_valid(monitor_1_io_in_a_valid),
		.io_in_a_bits_address(monitor_1_io_in_a_bits_address),
		.io_in_d_valid(monitor_1_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_1_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_1_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_1_io_in_d_bits_size),
		.io_in_d_bits_sink(monitor_1_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_1_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_1_io_in_d_bits_corrupt)
	);
	assign auto_in_1_a_ready = auto_out_a_ready & allowed_1;
	assign auto_in_1_d_valid = auto_out_d_valid & requestDOI_0_1;
	assign auto_in_1_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_1_d_bits_size = auto_out_d_bits_size;
	assign auto_in_1_d_bits_data = auto_out_d_bits_data;
	assign auto_in_1_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_in_0_a_ready = auto_out_a_ready & allowed_0;
	assign auto_in_0_d_valid = auto_out_d_valid & auto_out_d_bits_source;
	assign auto_in_0_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_0_d_bits_size = auto_out_d_bits_size;
	assign auto_in_0_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_0_d_bits_data = auto_out_d_bits_data;
	assign auto_out_a_valid = (idle ? _T_10 : _out_0_a_earlyValid_T_3);
	assign auto_out_a_bits_opcode = _T_45 | _T_46;
	assign auto_out_a_bits_param = (muxStateEarly_0 ? auto_in_0_a_bits_param : 3'h0);
	assign auto_out_a_bits_size = _T_39 | _T_40;
	assign auto_out_a_bits_source = (idle ? earlyWinner_0 : state_0);
	assign auto_out_a_bits_address = _T_33 | _T_34;
	assign auto_out_a_bits_mask = _T_30 | _T_31;
	assign auto_out_a_bits_data = (muxStateEarly_0 ? auto_in_0_a_bits_data : 32'h00000000);
	assign auto_out_d_ready = (auto_out_d_bits_source & auto_in_0_d_ready) | requestDOI_0_1;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_out_a_ready & allowed_0;
	assign monitor_io_in_a_valid = auto_in_0_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_0_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_0_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_0_a_bits_size;
	assign monitor_io_in_a_bits_address = auto_in_0_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_0_a_bits_mask;
	assign monitor_io_in_d_ready = auto_in_0_d_ready;
	assign monitor_io_in_d_valid = auto_out_d_valid & auto_out_d_bits_source;
	assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_io_in_d_bits_param = auto_out_d_bits_param;
	assign monitor_io_in_d_bits_size = auto_out_d_bits_size;
	assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink;
	assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied;
	assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign monitor_1_clock = clock;
	assign monitor_1_reset = reset;
	assign monitor_1_io_in_a_ready = auto_out_a_ready & allowed_1;
	assign monitor_1_io_in_a_valid = auto_in_1_a_valid;
	assign monitor_1_io_in_a_bits_address = auto_in_1_a_bits_address;
	assign monitor_1_io_in_d_valid = auto_out_d_valid & requestDOI_0_1;
	assign monitor_1_io_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign monitor_1_io_in_d_bits_param = auto_out_d_bits_param;
	assign monitor_1_io_in_d_bits_size = auto_out_d_bits_size;
	assign monitor_1_io_in_d_bits_sink = auto_out_d_bits_sink;
	assign monitor_1_io_in_d_bits_denied = auto_out_d_bits_denied;
	assign monitor_1_io_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	always @(posedge clock) begin
		if (reset)
			beatsLeft <= 10'h000;
		else if (latch) begin
			if (earlyWinner_0) begin
				if (beatsAI_opdata)
					beatsLeft <= beatsAI_decode;
				else
					beatsLeft <= 10'h000;
			end
			else
				beatsLeft <= 10'h000;
		end
		else
			beatsLeft <= _beatsLeft_T_4;
		if (reset)
			readys_mask <= 2'h3;
		else if (latch & |readys_valid)
			readys_mask <= _readys_mask_T_3;
		if (reset)
			state_0 <= 1'h0;
		else if (idle)
			state_0 <= earlyWinner_0;
		if (reset)
			state_1 <= 1'h0;
		else if (idle)
			state_1 <= earlyWinner_1;
	end
endmodule
module TLXbar_7 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module IntXbar_1 (
	auto_int_in_2_0,
	auto_int_in_1_0,
	auto_int_in_1_1,
	auto_int_in_0_0,
	auto_int_out_0,
	auto_int_out_1,
	auto_int_out_2,
	auto_int_out_3
);
	input auto_int_in_2_0;
	input auto_int_in_1_0;
	input auto_int_in_1_1;
	input auto_int_in_0_0;
	output wire auto_int_out_0;
	output wire auto_int_out_1;
	output wire auto_int_out_2;
	output wire auto_int_out_3;
	assign auto_int_out_0 = auto_int_in_0_0;
	assign auto_int_out_1 = auto_int_in_1_0;
	assign auto_int_out_2 = auto_int_in_1_1;
	assign auto_int_out_3 = auto_int_in_2_0;
endmodule
module BundleBridgeNexus_4 (
	auto_in,
	auto_out_0
);
	input auto_in;
	output wire auto_out_0;
	assign auto_out_0 = auto_in;
endmodule
module PMPChecker (
	io_prv,
	io_pmp_0_cfg_l,
	io_pmp_0_cfg_a,
	io_pmp_0_cfg_x,
	io_pmp_0_cfg_w,
	io_pmp_0_cfg_r,
	io_pmp_0_addr,
	io_pmp_0_mask,
	io_pmp_1_cfg_l,
	io_pmp_1_cfg_a,
	io_pmp_1_cfg_x,
	io_pmp_1_cfg_w,
	io_pmp_1_cfg_r,
	io_pmp_1_addr,
	io_pmp_1_mask,
	io_pmp_2_cfg_l,
	io_pmp_2_cfg_a,
	io_pmp_2_cfg_x,
	io_pmp_2_cfg_w,
	io_pmp_2_cfg_r,
	io_pmp_2_addr,
	io_pmp_2_mask,
	io_pmp_3_cfg_l,
	io_pmp_3_cfg_a,
	io_pmp_3_cfg_x,
	io_pmp_3_cfg_w,
	io_pmp_3_cfg_r,
	io_pmp_3_addr,
	io_pmp_3_mask,
	io_pmp_4_cfg_l,
	io_pmp_4_cfg_a,
	io_pmp_4_cfg_x,
	io_pmp_4_cfg_w,
	io_pmp_4_cfg_r,
	io_pmp_4_addr,
	io_pmp_4_mask,
	io_pmp_5_cfg_l,
	io_pmp_5_cfg_a,
	io_pmp_5_cfg_x,
	io_pmp_5_cfg_w,
	io_pmp_5_cfg_r,
	io_pmp_5_addr,
	io_pmp_5_mask,
	io_pmp_6_cfg_l,
	io_pmp_6_cfg_a,
	io_pmp_6_cfg_x,
	io_pmp_6_cfg_w,
	io_pmp_6_cfg_r,
	io_pmp_6_addr,
	io_pmp_6_mask,
	io_pmp_7_cfg_l,
	io_pmp_7_cfg_a,
	io_pmp_7_cfg_x,
	io_pmp_7_cfg_w,
	io_pmp_7_cfg_r,
	io_pmp_7_addr,
	io_pmp_7_mask,
	io_addr,
	io_r,
	io_w,
	io_x
);
	input [1:0] io_prv;
	input io_pmp_0_cfg_l;
	input [1:0] io_pmp_0_cfg_a;
	input io_pmp_0_cfg_x;
	input io_pmp_0_cfg_w;
	input io_pmp_0_cfg_r;
	input [29:0] io_pmp_0_addr;
	input [31:0] io_pmp_0_mask;
	input io_pmp_1_cfg_l;
	input [1:0] io_pmp_1_cfg_a;
	input io_pmp_1_cfg_x;
	input io_pmp_1_cfg_w;
	input io_pmp_1_cfg_r;
	input [29:0] io_pmp_1_addr;
	input [31:0] io_pmp_1_mask;
	input io_pmp_2_cfg_l;
	input [1:0] io_pmp_2_cfg_a;
	input io_pmp_2_cfg_x;
	input io_pmp_2_cfg_w;
	input io_pmp_2_cfg_r;
	input [29:0] io_pmp_2_addr;
	input [31:0] io_pmp_2_mask;
	input io_pmp_3_cfg_l;
	input [1:0] io_pmp_3_cfg_a;
	input io_pmp_3_cfg_x;
	input io_pmp_3_cfg_w;
	input io_pmp_3_cfg_r;
	input [29:0] io_pmp_3_addr;
	input [31:0] io_pmp_3_mask;
	input io_pmp_4_cfg_l;
	input [1:0] io_pmp_4_cfg_a;
	input io_pmp_4_cfg_x;
	input io_pmp_4_cfg_w;
	input io_pmp_4_cfg_r;
	input [29:0] io_pmp_4_addr;
	input [31:0] io_pmp_4_mask;
	input io_pmp_5_cfg_l;
	input [1:0] io_pmp_5_cfg_a;
	input io_pmp_5_cfg_x;
	input io_pmp_5_cfg_w;
	input io_pmp_5_cfg_r;
	input [29:0] io_pmp_5_addr;
	input [31:0] io_pmp_5_mask;
	input io_pmp_6_cfg_l;
	input [1:0] io_pmp_6_cfg_a;
	input io_pmp_6_cfg_x;
	input io_pmp_6_cfg_w;
	input io_pmp_6_cfg_r;
	input [29:0] io_pmp_6_addr;
	input [31:0] io_pmp_6_mask;
	input io_pmp_7_cfg_l;
	input [1:0] io_pmp_7_cfg_a;
	input io_pmp_7_cfg_x;
	input io_pmp_7_cfg_w;
	input io_pmp_7_cfg_r;
	input [29:0] io_pmp_7_addr;
	input [31:0] io_pmp_7_mask;
	input [31:0] io_addr;
	output wire io_r;
	output wire io_w;
	output wire io_x;
	wire default_ = io_prv > 2'h1;
	wire [31:0] _res_hit_T_1 = {io_pmp_7_addr, 2'h0};
	wire [31:0] _res_hit_T_2 = ~_res_hit_T_1;
	wire [31:0] _res_hit_T_3 = _res_hit_T_2 | 32'h00000003;
	wire [31:0] _res_hit_T_4 = ~_res_hit_T_3;
	wire [31:0] _res_hit_T_5 = io_addr ^ _res_hit_T_4;
	wire [31:0] _res_hit_T_6 = ~io_pmp_7_mask;
	wire [31:0] _res_hit_T_7 = _res_hit_T_5 & _res_hit_T_6;
	wire _res_hit_T_8 = _res_hit_T_7 == 32'h00000000;
	wire [31:0] _res_hit_T_14 = {io_pmp_6_addr, 2'h0};
	wire [31:0] _res_hit_T_15 = ~_res_hit_T_14;
	wire [31:0] _res_hit_T_16 = _res_hit_T_15 | 32'h00000003;
	wire [31:0] _res_hit_T_17 = ~_res_hit_T_16;
	wire _res_hit_T_18 = io_addr < _res_hit_T_17;
	wire _res_hit_T_19 = ~_res_hit_T_18;
	wire _res_hit_T_24 = io_addr < _res_hit_T_4;
	wire _res_hit_T_25 = _res_hit_T_19 & _res_hit_T_24;
	wire res_hit = (io_pmp_7_cfg_a[1] ? _res_hit_T_8 : io_pmp_7_cfg_a[0] & _res_hit_T_25);
	wire res_ignore = default_ & ~io_pmp_7_cfg_l;
	wire res_cur_cfg_r = io_pmp_7_cfg_r | res_ignore;
	wire res_cur_cfg_w = io_pmp_7_cfg_w | res_ignore;
	wire res_cur_cfg_x = io_pmp_7_cfg_x | res_ignore;
	wire _res_T_44_cfg_x = (res_hit ? res_cur_cfg_x : default_);
	wire _res_T_44_cfg_w = (res_hit ? res_cur_cfg_w : default_);
	wire _res_T_44_cfg_r = (res_hit ? res_cur_cfg_r : default_);
	wire [31:0] _res_hit_T_32 = io_addr ^ _res_hit_T_17;
	wire [31:0] _res_hit_T_33 = ~io_pmp_6_mask;
	wire [31:0] _res_hit_T_34 = _res_hit_T_32 & _res_hit_T_33;
	wire _res_hit_T_35 = _res_hit_T_34 == 32'h00000000;
	wire [31:0] _res_hit_T_41 = {io_pmp_5_addr, 2'h0};
	wire [31:0] _res_hit_T_42 = ~_res_hit_T_41;
	wire [31:0] _res_hit_T_43 = _res_hit_T_42 | 32'h00000003;
	wire [31:0] _res_hit_T_44 = ~_res_hit_T_43;
	wire _res_hit_T_45 = io_addr < _res_hit_T_44;
	wire _res_hit_T_46 = ~_res_hit_T_45;
	wire _res_hit_T_52 = _res_hit_T_46 & _res_hit_T_18;
	wire res_hit_1 = (io_pmp_6_cfg_a[1] ? _res_hit_T_35 : io_pmp_6_cfg_a[0] & _res_hit_T_52);
	wire res_ignore_1 = default_ & ~io_pmp_6_cfg_l;
	wire res_cur_1_cfg_r = io_pmp_6_cfg_r | res_ignore_1;
	wire res_cur_1_cfg_w = io_pmp_6_cfg_w | res_ignore_1;
	wire res_cur_1_cfg_x = io_pmp_6_cfg_x | res_ignore_1;
	wire _res_T_89_cfg_x = (res_hit_1 ? res_cur_1_cfg_x : _res_T_44_cfg_x);
	wire _res_T_89_cfg_w = (res_hit_1 ? res_cur_1_cfg_w : _res_T_44_cfg_w);
	wire _res_T_89_cfg_r = (res_hit_1 ? res_cur_1_cfg_r : _res_T_44_cfg_r);
	wire [31:0] _res_hit_T_59 = io_addr ^ _res_hit_T_44;
	wire [31:0] _res_hit_T_60 = ~io_pmp_5_mask;
	wire [31:0] _res_hit_T_61 = _res_hit_T_59 & _res_hit_T_60;
	wire _res_hit_T_62 = _res_hit_T_61 == 32'h00000000;
	wire [31:0] _res_hit_T_68 = {io_pmp_4_addr, 2'h0};
	wire [31:0] _res_hit_T_69 = ~_res_hit_T_68;
	wire [31:0] _res_hit_T_70 = _res_hit_T_69 | 32'h00000003;
	wire [31:0] _res_hit_T_71 = ~_res_hit_T_70;
	wire _res_hit_T_72 = io_addr < _res_hit_T_71;
	wire _res_hit_T_73 = ~_res_hit_T_72;
	wire _res_hit_T_79 = _res_hit_T_73 & _res_hit_T_45;
	wire res_hit_2 = (io_pmp_5_cfg_a[1] ? _res_hit_T_62 : io_pmp_5_cfg_a[0] & _res_hit_T_79);
	wire res_ignore_2 = default_ & ~io_pmp_5_cfg_l;
	wire res_cur_2_cfg_r = io_pmp_5_cfg_r | res_ignore_2;
	wire res_cur_2_cfg_w = io_pmp_5_cfg_w | res_ignore_2;
	wire res_cur_2_cfg_x = io_pmp_5_cfg_x | res_ignore_2;
	wire _res_T_134_cfg_x = (res_hit_2 ? res_cur_2_cfg_x : _res_T_89_cfg_x);
	wire _res_T_134_cfg_w = (res_hit_2 ? res_cur_2_cfg_w : _res_T_89_cfg_w);
	wire _res_T_134_cfg_r = (res_hit_2 ? res_cur_2_cfg_r : _res_T_89_cfg_r);
	wire [31:0] _res_hit_T_86 = io_addr ^ _res_hit_T_71;
	wire [31:0] _res_hit_T_87 = ~io_pmp_4_mask;
	wire [31:0] _res_hit_T_88 = _res_hit_T_86 & _res_hit_T_87;
	wire _res_hit_T_89 = _res_hit_T_88 == 32'h00000000;
	wire [31:0] _res_hit_T_95 = {io_pmp_3_addr, 2'h0};
	wire [31:0] _res_hit_T_96 = ~_res_hit_T_95;
	wire [31:0] _res_hit_T_97 = _res_hit_T_96 | 32'h00000003;
	wire [31:0] _res_hit_T_98 = ~_res_hit_T_97;
	wire _res_hit_T_99 = io_addr < _res_hit_T_98;
	wire _res_hit_T_100 = ~_res_hit_T_99;
	wire _res_hit_T_106 = _res_hit_T_100 & _res_hit_T_72;
	wire res_hit_3 = (io_pmp_4_cfg_a[1] ? _res_hit_T_89 : io_pmp_4_cfg_a[0] & _res_hit_T_106);
	wire res_ignore_3 = default_ & ~io_pmp_4_cfg_l;
	wire res_cur_3_cfg_r = io_pmp_4_cfg_r | res_ignore_3;
	wire res_cur_3_cfg_w = io_pmp_4_cfg_w | res_ignore_3;
	wire res_cur_3_cfg_x = io_pmp_4_cfg_x | res_ignore_3;
	wire _res_T_179_cfg_x = (res_hit_3 ? res_cur_3_cfg_x : _res_T_134_cfg_x);
	wire _res_T_179_cfg_w = (res_hit_3 ? res_cur_3_cfg_w : _res_T_134_cfg_w);
	wire _res_T_179_cfg_r = (res_hit_3 ? res_cur_3_cfg_r : _res_T_134_cfg_r);
	wire [31:0] _res_hit_T_113 = io_addr ^ _res_hit_T_98;
	wire [31:0] _res_hit_T_114 = ~io_pmp_3_mask;
	wire [31:0] _res_hit_T_115 = _res_hit_T_113 & _res_hit_T_114;
	wire _res_hit_T_116 = _res_hit_T_115 == 32'h00000000;
	wire [31:0] _res_hit_T_122 = {io_pmp_2_addr, 2'h0};
	wire [31:0] _res_hit_T_123 = ~_res_hit_T_122;
	wire [31:0] _res_hit_T_124 = _res_hit_T_123 | 32'h00000003;
	wire [31:0] _res_hit_T_125 = ~_res_hit_T_124;
	wire _res_hit_T_126 = io_addr < _res_hit_T_125;
	wire _res_hit_T_127 = ~_res_hit_T_126;
	wire _res_hit_T_133 = _res_hit_T_127 & _res_hit_T_99;
	wire res_hit_4 = (io_pmp_3_cfg_a[1] ? _res_hit_T_116 : io_pmp_3_cfg_a[0] & _res_hit_T_133);
	wire res_ignore_4 = default_ & ~io_pmp_3_cfg_l;
	wire res_cur_4_cfg_r = io_pmp_3_cfg_r | res_ignore_4;
	wire res_cur_4_cfg_w = io_pmp_3_cfg_w | res_ignore_4;
	wire res_cur_4_cfg_x = io_pmp_3_cfg_x | res_ignore_4;
	wire _res_T_224_cfg_x = (res_hit_4 ? res_cur_4_cfg_x : _res_T_179_cfg_x);
	wire _res_T_224_cfg_w = (res_hit_4 ? res_cur_4_cfg_w : _res_T_179_cfg_w);
	wire _res_T_224_cfg_r = (res_hit_4 ? res_cur_4_cfg_r : _res_T_179_cfg_r);
	wire [31:0] _res_hit_T_140 = io_addr ^ _res_hit_T_125;
	wire [31:0] _res_hit_T_141 = ~io_pmp_2_mask;
	wire [31:0] _res_hit_T_142 = _res_hit_T_140 & _res_hit_T_141;
	wire _res_hit_T_143 = _res_hit_T_142 == 32'h00000000;
	wire [31:0] _res_hit_T_149 = {io_pmp_1_addr, 2'h0};
	wire [31:0] _res_hit_T_150 = ~_res_hit_T_149;
	wire [31:0] _res_hit_T_151 = _res_hit_T_150 | 32'h00000003;
	wire [31:0] _res_hit_T_152 = ~_res_hit_T_151;
	wire _res_hit_T_153 = io_addr < _res_hit_T_152;
	wire _res_hit_T_154 = ~_res_hit_T_153;
	wire _res_hit_T_160 = _res_hit_T_154 & _res_hit_T_126;
	wire res_hit_5 = (io_pmp_2_cfg_a[1] ? _res_hit_T_143 : io_pmp_2_cfg_a[0] & _res_hit_T_160);
	wire res_ignore_5 = default_ & ~io_pmp_2_cfg_l;
	wire res_cur_5_cfg_r = io_pmp_2_cfg_r | res_ignore_5;
	wire res_cur_5_cfg_w = io_pmp_2_cfg_w | res_ignore_5;
	wire res_cur_5_cfg_x = io_pmp_2_cfg_x | res_ignore_5;
	wire _res_T_269_cfg_x = (res_hit_5 ? res_cur_5_cfg_x : _res_T_224_cfg_x);
	wire _res_T_269_cfg_w = (res_hit_5 ? res_cur_5_cfg_w : _res_T_224_cfg_w);
	wire _res_T_269_cfg_r = (res_hit_5 ? res_cur_5_cfg_r : _res_T_224_cfg_r);
	wire [31:0] _res_hit_T_167 = io_addr ^ _res_hit_T_152;
	wire [31:0] _res_hit_T_168 = ~io_pmp_1_mask;
	wire [31:0] _res_hit_T_169 = _res_hit_T_167 & _res_hit_T_168;
	wire _res_hit_T_170 = _res_hit_T_169 == 32'h00000000;
	wire [31:0] _res_hit_T_176 = {io_pmp_0_addr, 2'h0};
	wire [31:0] _res_hit_T_177 = ~_res_hit_T_176;
	wire [31:0] _res_hit_T_178 = _res_hit_T_177 | 32'h00000003;
	wire [31:0] _res_hit_T_179 = ~_res_hit_T_178;
	wire _res_hit_T_180 = io_addr < _res_hit_T_179;
	wire _res_hit_T_181 = ~_res_hit_T_180;
	wire _res_hit_T_187 = _res_hit_T_181 & _res_hit_T_153;
	wire res_hit_6 = (io_pmp_1_cfg_a[1] ? _res_hit_T_170 : io_pmp_1_cfg_a[0] & _res_hit_T_187);
	wire res_ignore_6 = default_ & ~io_pmp_1_cfg_l;
	wire res_cur_6_cfg_r = io_pmp_1_cfg_r | res_ignore_6;
	wire res_cur_6_cfg_w = io_pmp_1_cfg_w | res_ignore_6;
	wire res_cur_6_cfg_x = io_pmp_1_cfg_x | res_ignore_6;
	wire _res_T_314_cfg_x = (res_hit_6 ? res_cur_6_cfg_x : _res_T_269_cfg_x);
	wire _res_T_314_cfg_w = (res_hit_6 ? res_cur_6_cfg_w : _res_T_269_cfg_w);
	wire _res_T_314_cfg_r = (res_hit_6 ? res_cur_6_cfg_r : _res_T_269_cfg_r);
	wire [31:0] _res_hit_T_194 = io_addr ^ _res_hit_T_179;
	wire [31:0] _res_hit_T_195 = ~io_pmp_0_mask;
	wire [31:0] _res_hit_T_196 = _res_hit_T_194 & _res_hit_T_195;
	wire _res_hit_T_197 = _res_hit_T_196 == 32'h00000000;
	wire res_hit_7 = (io_pmp_0_cfg_a[1] ? _res_hit_T_197 : io_pmp_0_cfg_a[0] & _res_hit_T_180);
	wire res_ignore_7 = default_ & ~io_pmp_0_cfg_l;
	wire res_cur_7_cfg_r = io_pmp_0_cfg_r | res_ignore_7;
	wire res_cur_7_cfg_w = io_pmp_0_cfg_w | res_ignore_7;
	wire res_cur_7_cfg_x = io_pmp_0_cfg_x | res_ignore_7;
	assign io_r = (res_hit_7 ? res_cur_7_cfg_r : _res_T_314_cfg_r);
	assign io_w = (res_hit_7 ? res_cur_7_cfg_w : _res_T_314_cfg_w);
	assign io_x = (res_hit_7 ? res_cur_7_cfg_x : _res_T_314_cfg_x);
endmodule
module TLB (
	io_req_valid,
	io_req_bits_vaddr,
	io_req_bits_size,
	io_req_bits_cmd,
	io_req_bits_prv,
	io_resp_paddr,
	io_resp_pf_ld,
	io_resp_pf_st,
	io_resp_ae_ld,
	io_resp_ae_st,
	io_resp_ma_ld,
	io_resp_ma_st,
	io_ptw_status_debug,
	io_ptw_pmp_0_cfg_l,
	io_ptw_pmp_0_cfg_a,
	io_ptw_pmp_0_cfg_x,
	io_ptw_pmp_0_cfg_w,
	io_ptw_pmp_0_cfg_r,
	io_ptw_pmp_0_addr,
	io_ptw_pmp_0_mask,
	io_ptw_pmp_1_cfg_l,
	io_ptw_pmp_1_cfg_a,
	io_ptw_pmp_1_cfg_x,
	io_ptw_pmp_1_cfg_w,
	io_ptw_pmp_1_cfg_r,
	io_ptw_pmp_1_addr,
	io_ptw_pmp_1_mask,
	io_ptw_pmp_2_cfg_l,
	io_ptw_pmp_2_cfg_a,
	io_ptw_pmp_2_cfg_x,
	io_ptw_pmp_2_cfg_w,
	io_ptw_pmp_2_cfg_r,
	io_ptw_pmp_2_addr,
	io_ptw_pmp_2_mask,
	io_ptw_pmp_3_cfg_l,
	io_ptw_pmp_3_cfg_a,
	io_ptw_pmp_3_cfg_x,
	io_ptw_pmp_3_cfg_w,
	io_ptw_pmp_3_cfg_r,
	io_ptw_pmp_3_addr,
	io_ptw_pmp_3_mask,
	io_ptw_pmp_4_cfg_l,
	io_ptw_pmp_4_cfg_a,
	io_ptw_pmp_4_cfg_x,
	io_ptw_pmp_4_cfg_w,
	io_ptw_pmp_4_cfg_r,
	io_ptw_pmp_4_addr,
	io_ptw_pmp_4_mask,
	io_ptw_pmp_5_cfg_l,
	io_ptw_pmp_5_cfg_a,
	io_ptw_pmp_5_cfg_x,
	io_ptw_pmp_5_cfg_w,
	io_ptw_pmp_5_cfg_r,
	io_ptw_pmp_5_addr,
	io_ptw_pmp_5_mask,
	io_ptw_pmp_6_cfg_l,
	io_ptw_pmp_6_cfg_a,
	io_ptw_pmp_6_cfg_x,
	io_ptw_pmp_6_cfg_w,
	io_ptw_pmp_6_cfg_r,
	io_ptw_pmp_6_addr,
	io_ptw_pmp_6_mask,
	io_ptw_pmp_7_cfg_l,
	io_ptw_pmp_7_cfg_a,
	io_ptw_pmp_7_cfg_x,
	io_ptw_pmp_7_cfg_w,
	io_ptw_pmp_7_cfg_r,
	io_ptw_pmp_7_addr,
	io_ptw_pmp_7_mask
);
	input io_req_valid;
	input [31:0] io_req_bits_vaddr;
	input [1:0] io_req_bits_size;
	input [4:0] io_req_bits_cmd;
	input [1:0] io_req_bits_prv;
	output wire [31:0] io_resp_paddr;
	output wire io_resp_pf_ld;
	output wire io_resp_pf_st;
	output wire io_resp_ae_ld;
	output wire io_resp_ae_st;
	output wire io_resp_ma_ld;
	output wire io_resp_ma_st;
	input io_ptw_status_debug;
	input io_ptw_pmp_0_cfg_l;
	input [1:0] io_ptw_pmp_0_cfg_a;
	input io_ptw_pmp_0_cfg_x;
	input io_ptw_pmp_0_cfg_w;
	input io_ptw_pmp_0_cfg_r;
	input [29:0] io_ptw_pmp_0_addr;
	input [31:0] io_ptw_pmp_0_mask;
	input io_ptw_pmp_1_cfg_l;
	input [1:0] io_ptw_pmp_1_cfg_a;
	input io_ptw_pmp_1_cfg_x;
	input io_ptw_pmp_1_cfg_w;
	input io_ptw_pmp_1_cfg_r;
	input [29:0] io_ptw_pmp_1_addr;
	input [31:0] io_ptw_pmp_1_mask;
	input io_ptw_pmp_2_cfg_l;
	input [1:0] io_ptw_pmp_2_cfg_a;
	input io_ptw_pmp_2_cfg_x;
	input io_ptw_pmp_2_cfg_w;
	input io_ptw_pmp_2_cfg_r;
	input [29:0] io_ptw_pmp_2_addr;
	input [31:0] io_ptw_pmp_2_mask;
	input io_ptw_pmp_3_cfg_l;
	input [1:0] io_ptw_pmp_3_cfg_a;
	input io_ptw_pmp_3_cfg_x;
	input io_ptw_pmp_3_cfg_w;
	input io_ptw_pmp_3_cfg_r;
	input [29:0] io_ptw_pmp_3_addr;
	input [31:0] io_ptw_pmp_3_mask;
	input io_ptw_pmp_4_cfg_l;
	input [1:0] io_ptw_pmp_4_cfg_a;
	input io_ptw_pmp_4_cfg_x;
	input io_ptw_pmp_4_cfg_w;
	input io_ptw_pmp_4_cfg_r;
	input [29:0] io_ptw_pmp_4_addr;
	input [31:0] io_ptw_pmp_4_mask;
	input io_ptw_pmp_5_cfg_l;
	input [1:0] io_ptw_pmp_5_cfg_a;
	input io_ptw_pmp_5_cfg_x;
	input io_ptw_pmp_5_cfg_w;
	input io_ptw_pmp_5_cfg_r;
	input [29:0] io_ptw_pmp_5_addr;
	input [31:0] io_ptw_pmp_5_mask;
	input io_ptw_pmp_6_cfg_l;
	input [1:0] io_ptw_pmp_6_cfg_a;
	input io_ptw_pmp_6_cfg_x;
	input io_ptw_pmp_6_cfg_w;
	input io_ptw_pmp_6_cfg_r;
	input [29:0] io_ptw_pmp_6_addr;
	input [31:0] io_ptw_pmp_6_mask;
	input io_ptw_pmp_7_cfg_l;
	input [1:0] io_ptw_pmp_7_cfg_a;
	input io_ptw_pmp_7_cfg_x;
	input io_ptw_pmp_7_cfg_w;
	input io_ptw_pmp_7_cfg_r;
	input [29:0] io_ptw_pmp_7_addr;
	input [31:0] io_ptw_pmp_7_mask;
	wire [1:0] pmp_io_prv;
	wire pmp_io_pmp_0_cfg_l;
	wire [1:0] pmp_io_pmp_0_cfg_a;
	wire pmp_io_pmp_0_cfg_x;
	wire pmp_io_pmp_0_cfg_w;
	wire pmp_io_pmp_0_cfg_r;
	wire [29:0] pmp_io_pmp_0_addr;
	wire [31:0] pmp_io_pmp_0_mask;
	wire pmp_io_pmp_1_cfg_l;
	wire [1:0] pmp_io_pmp_1_cfg_a;
	wire pmp_io_pmp_1_cfg_x;
	wire pmp_io_pmp_1_cfg_w;
	wire pmp_io_pmp_1_cfg_r;
	wire [29:0] pmp_io_pmp_1_addr;
	wire [31:0] pmp_io_pmp_1_mask;
	wire pmp_io_pmp_2_cfg_l;
	wire [1:0] pmp_io_pmp_2_cfg_a;
	wire pmp_io_pmp_2_cfg_x;
	wire pmp_io_pmp_2_cfg_w;
	wire pmp_io_pmp_2_cfg_r;
	wire [29:0] pmp_io_pmp_2_addr;
	wire [31:0] pmp_io_pmp_2_mask;
	wire pmp_io_pmp_3_cfg_l;
	wire [1:0] pmp_io_pmp_3_cfg_a;
	wire pmp_io_pmp_3_cfg_x;
	wire pmp_io_pmp_3_cfg_w;
	wire pmp_io_pmp_3_cfg_r;
	wire [29:0] pmp_io_pmp_3_addr;
	wire [31:0] pmp_io_pmp_3_mask;
	wire pmp_io_pmp_4_cfg_l;
	wire [1:0] pmp_io_pmp_4_cfg_a;
	wire pmp_io_pmp_4_cfg_x;
	wire pmp_io_pmp_4_cfg_w;
	wire pmp_io_pmp_4_cfg_r;
	wire [29:0] pmp_io_pmp_4_addr;
	wire [31:0] pmp_io_pmp_4_mask;
	wire pmp_io_pmp_5_cfg_l;
	wire [1:0] pmp_io_pmp_5_cfg_a;
	wire pmp_io_pmp_5_cfg_x;
	wire pmp_io_pmp_5_cfg_w;
	wire pmp_io_pmp_5_cfg_r;
	wire [29:0] pmp_io_pmp_5_addr;
	wire [31:0] pmp_io_pmp_5_mask;
	wire pmp_io_pmp_6_cfg_l;
	wire [1:0] pmp_io_pmp_6_cfg_a;
	wire pmp_io_pmp_6_cfg_x;
	wire pmp_io_pmp_6_cfg_w;
	wire pmp_io_pmp_6_cfg_r;
	wire [29:0] pmp_io_pmp_6_addr;
	wire [31:0] pmp_io_pmp_6_mask;
	wire pmp_io_pmp_7_cfg_l;
	wire [1:0] pmp_io_pmp_7_cfg_a;
	wire pmp_io_pmp_7_cfg_x;
	wire pmp_io_pmp_7_cfg_w;
	wire pmp_io_pmp_7_cfg_r;
	wire [29:0] pmp_io_pmp_7_addr;
	wire [31:0] pmp_io_pmp_7_mask;
	wire [31:0] pmp_io_addr;
	wire pmp_io_r;
	wire pmp_io_w;
	wire pmp_io_x;
	wire [19:0] vpn = io_req_bits_vaddr[31:12];
	wire [19:0] mpu_ppn = io_req_bits_vaddr[31:12];
	wire [31:0] mpu_physaddr = {mpu_ppn, io_req_bits_vaddr[11:0]};
	wire [2:0] mpu_priv = {io_ptw_status_debug, io_req_bits_prv};
	wire [31:0] _legal_address_T = mpu_physaddr ^ 32'h00003000;
	wire [32:0] _legal_address_T_1 = {1'b0, $signed(_legal_address_T)};
	wire [32:0] _legal_address_T_3 = $signed(_legal_address_T_1) & -33'sh000001000;
	wire _legal_address_T_4 = $signed(_legal_address_T_3) == 33'sh000000000;
	wire [31:0] _legal_address_T_5 = mpu_physaddr ^ 32'h00004000;
	wire [32:0] _legal_address_T_6 = {1'b0, $signed(_legal_address_T_5)};
	wire [32:0] _legal_address_T_8 = $signed(_legal_address_T_6) & -33'sh000001000;
	wire _legal_address_T_9 = $signed(_legal_address_T_8) == 33'sh000000000;
	wire [31:0] _legal_address_T_10 = mpu_physaddr ^ 32'h10000000;
	wire [32:0] _legal_address_T_11 = {1'b0, $signed(_legal_address_T_10)};
	wire [32:0] _legal_address_T_13 = $signed(_legal_address_T_11) & -33'sh000001000;
	wire _legal_address_T_14 = $signed(_legal_address_T_13) == 33'sh000000000;
	wire [31:0] _legal_address_T_15 = mpu_physaddr ^ 32'h00020000;
	wire [32:0] _legal_address_T_16 = {1'b0, $signed(_legal_address_T_15)};
	wire [32:0] _legal_address_T_18 = $signed(_legal_address_T_16) & -33'sh000010000;
	wire _legal_address_T_19 = $signed(_legal_address_T_18) == 33'sh000000000;
	wire [31:0] _legal_address_T_20 = mpu_physaddr ^ 32'h54000000;
	wire [32:0] _legal_address_T_21 = {1'b0, $signed(_legal_address_T_20)};
	wire [32:0] _legal_address_T_23 = $signed(_legal_address_T_21) & -33'sh000001000;
	wire _legal_address_T_24 = $signed(_legal_address_T_23) == 33'sh000000000;
	wire [31:0] _legal_address_T_25 = mpu_physaddr ^ 32'h0c000000;
	wire [32:0] _legal_address_T_26 = {1'b0, $signed(_legal_address_T_25)};
	wire [32:0] _legal_address_T_28 = $signed(_legal_address_T_26) & -33'sh004000000;
	wire _legal_address_T_29 = $signed(_legal_address_T_28) == 33'sh000000000;
	wire [31:0] _legal_address_T_30 = mpu_physaddr ^ 32'h02000000;
	wire [32:0] _legal_address_T_31 = {1'b0, $signed(_legal_address_T_30)};
	wire [32:0] _legal_address_T_33 = $signed(_legal_address_T_31) & -33'sh000010000;
	wire _legal_address_T_34 = $signed(_legal_address_T_33) == 33'sh000000000;
	wire [32:0] _legal_address_T_36 = {1'b0, $signed(mpu_physaddr)};
	wire [32:0] _legal_address_T_38 = $signed(_legal_address_T_36) & -33'sh000001000;
	wire _legal_address_T_39 = $signed(_legal_address_T_38) == 33'sh000000000;
	wire [31:0] _legal_address_T_40 = mpu_physaddr ^ 32'h80000000;
	wire [32:0] _legal_address_T_41 = {1'b0, $signed(_legal_address_T_40)};
	wire [32:0] _legal_address_T_43 = $signed(_legal_address_T_41) & -33'sh000004000;
	wire _legal_address_T_44 = $signed(_legal_address_T_43) == 33'sh000000000;
	wire [31:0] _legal_address_T_45 = mpu_physaddr ^ 32'h00010000;
	wire [32:0] _legal_address_T_46 = {1'b0, $signed(_legal_address_T_45)};
	wire [32:0] _legal_address_T_48 = $signed(_legal_address_T_46) & -33'sh000010000;
	wire _legal_address_T_49 = $signed(_legal_address_T_48) == 33'sh000000000;
	wire [31:0] _legal_address_T_50 = mpu_physaddr ^ 32'h00100000;
	wire [32:0] _legal_address_T_51 = {1'b0, $signed(_legal_address_T_50)};
	wire [32:0] _legal_address_T_53 = $signed(_legal_address_T_51) & -33'sh000001000;
	wire _legal_address_T_54 = $signed(_legal_address_T_53) == 33'sh000000000;
	wire [31:0] _legal_address_T_55 = mpu_physaddr ^ 32'h00110000;
	wire [32:0] _legal_address_T_56 = {1'b0, $signed(_legal_address_T_55)};
	wire [32:0] _legal_address_T_58 = $signed(_legal_address_T_56) & -33'sh000001000;
	wire _legal_address_T_59 = $signed(_legal_address_T_58) == 33'sh000000000;
	wire legal_address = ((((((((((_legal_address_T_4 | _legal_address_T_9) | _legal_address_T_14) | _legal_address_T_19) | _legal_address_T_24) | _legal_address_T_29) | _legal_address_T_34) | _legal_address_T_39) | _legal_address_T_44) | _legal_address_T_49) | _legal_address_T_54) | _legal_address_T_59;
	wire deny_access_to_debug = (mpu_priv <= 3'h3) & _legal_address_T_39;
	wire _prot_r_T_6 = ~deny_access_to_debug;
	wire prot_r = (legal_address & ~deny_access_to_debug) & pmp_io_r;
	wire [32:0] _prot_w_T_3 = $signed(_legal_address_T_36) & 33'sh098130000;
	wire _prot_w_T_4 = $signed(_prot_w_T_3) == 33'sh000000000;
	wire [32:0] _prot_w_T_8 = $signed(_legal_address_T_51) & 33'sh09a120000;
	wire _prot_w_T_9 = $signed(_prot_w_T_8) == 33'sh000000000;
	wire [31:0] _prot_w_T_10 = mpu_physaddr ^ 32'h08000000;
	wire [32:0] _prot_w_T_11 = {1'b0, $signed(_prot_w_T_10)};
	wire [32:0] _prot_w_T_13 = $signed(_prot_w_T_11) & 33'sh098000000;
	wire _prot_w_T_14 = $signed(_prot_w_T_13) == 33'sh000000000;
	wire [32:0] _prot_w_T_18 = $signed(_legal_address_T_11) & 33'sh09a130000;
	wire _prot_w_T_19 = $signed(_prot_w_T_18) == 33'sh000000000;
	wire [32:0] _prot_w_T_23 = $signed(_legal_address_T_41) & 33'sh09a130000;
	wire _prot_w_T_24 = $signed(_prot_w_T_23) == 33'sh000000000;
	wire _prot_w_T_28 = (((_prot_w_T_4 | _prot_w_T_9) | _prot_w_T_14) | _prot_w_T_19) | _prot_w_T_24;
	wire _prot_w_T_43 = legal_address & _prot_w_T_28;
	wire prot_w = (_prot_w_T_43 & _prot_r_T_6) & pmp_io_w;
	wire [32:0] _prot_x_T_36 = $signed(_legal_address_T_31) & 33'sh096130000;
	wire _prot_x_T_37 = $signed(_prot_x_T_36) == 33'sh000000000;
	wire [31:0] _prot_x_T_38 = mpu_physaddr ^ 32'h04000000;
	wire [32:0] _prot_x_T_39 = {1'b0, $signed(_prot_x_T_38)};
	wire [32:0] _prot_x_T_41 = $signed(_prot_x_T_39) & 33'sh094000000;
	wire _prot_x_T_42 = $signed(_prot_x_T_41) == 33'sh000000000;
	wire [31:0] _prot_x_T_43 = mpu_physaddr ^ 32'h14000000;
	wire [32:0] _prot_x_T_44 = {1'b0, $signed(_prot_x_T_43)};
	wire [32:0] _prot_eff_T_32 = $signed(_legal_address_T_36) & 33'sh096132000;
	wire _prot_eff_T_33 = $signed(_prot_eff_T_32) == 33'sh000000000;
	wire [32:0] _prot_eff_T_37 = $signed(_legal_address_T_51) & 33'sh096122000;
	wire _prot_eff_T_38 = $signed(_prot_eff_T_37) == 33'sh000000000;
	wire [32:0] _prot_eff_T_52 = $signed(_prot_x_T_44) & 33'sh096132000;
	wire _prot_eff_T_53 = $signed(_prot_eff_T_52) == 33'sh000000000;
	wire _prot_eff_T_57 = (((_prot_eff_T_33 | _prot_eff_T_38) | _prot_x_T_37) | _prot_x_T_42) | _prot_eff_T_53;
	wire prot_eff = legal_address & _prot_eff_T_57;
	wire [1:0] _pr_array_T_1 = (prot_r ? 2'h3 : 2'h0);
	wire [6:0] pr_array = {_pr_array_T_1, 5'h00};
	wire [1:0] _pw_array_T_1 = (prot_w ? 2'h3 : 2'h0);
	wire [6:0] pw_array = {_pw_array_T_1, 5'h00};
	wire [1:0] _eff_array_T_1 = (prot_eff ? 2'h3 : 2'h0);
	wire [6:0] eff_array = {_eff_array_T_1, 5'h00};
	wire [1:0] _ppp_array_T_1 = (_prot_w_T_43 ? 2'h3 : 2'h0);
	wire [6:0] ppp_array = {_ppp_array_T_1, 5'h00};
	wire [3:0] _misaligned_T = 4'h1 << io_req_bits_size;
	wire [3:0] _misaligned_T_2 = _misaligned_T - 4'h1;
	wire [31:0] _GEN_144 = {28'd0, _misaligned_T_2};
	wire [31:0] _misaligned_T_3 = io_req_bits_vaddr & _GEN_144;
	wire misaligned = |_misaligned_T_3;
	wire _cmd_lrsc_T = io_req_bits_cmd == 5'h06;
	wire _cmd_lrsc_T_1 = io_req_bits_cmd == 5'h07;
	wire cmd_lrsc = _cmd_lrsc_T | _cmd_lrsc_T_1;
	wire _cmd_amo_logical_T = io_req_bits_cmd == 5'h04;
	wire _cmd_amo_logical_T_1 = io_req_bits_cmd == 5'h09;
	wire _cmd_amo_logical_T_2 = io_req_bits_cmd == 5'h0a;
	wire _cmd_amo_logical_T_3 = io_req_bits_cmd == 5'h0b;
	wire cmd_amo_logical = ((_cmd_amo_logical_T | _cmd_amo_logical_T_1) | _cmd_amo_logical_T_2) | _cmd_amo_logical_T_3;
	wire _cmd_amo_arithmetic_T = io_req_bits_cmd == 5'h08;
	wire _cmd_amo_arithmetic_T_1 = io_req_bits_cmd == 5'h0c;
	wire _cmd_amo_arithmetic_T_2 = io_req_bits_cmd == 5'h0d;
	wire _cmd_amo_arithmetic_T_3 = io_req_bits_cmd == 5'h0e;
	wire _cmd_amo_arithmetic_T_4 = io_req_bits_cmd == 5'h0f;
	wire cmd_amo_arithmetic = (((_cmd_amo_arithmetic_T | _cmd_amo_arithmetic_T_1) | _cmd_amo_arithmetic_T_2) | _cmd_amo_arithmetic_T_3) | _cmd_amo_arithmetic_T_4;
	wire cmd_put_partial = io_req_bits_cmd == 5'h11;
	wire _cmd_read_T = io_req_bits_cmd == 5'h00;
	wire _cmd_read_T_1 = io_req_bits_cmd == 5'h10;
	wire _cmd_read_T_6 = ((_cmd_read_T | _cmd_read_T_1) | _cmd_lrsc_T) | _cmd_lrsc_T_1;
	wire _cmd_read_T_23 = cmd_amo_logical | cmd_amo_arithmetic;
	wire cmd_read = _cmd_read_T_6 | _cmd_read_T_23;
	wire cmd_write = (((io_req_bits_cmd == 5'h01) | cmd_put_partial) | _cmd_lrsc_T_1) | _cmd_read_T_23;
	wire _cmd_write_perms_T = io_req_bits_cmd == 5'h05;
	wire _cmd_write_perms_T_1 = io_req_bits_cmd == 5'h17;
	wire _cmd_write_perms_T_2 = _cmd_write_perms_T | _cmd_write_perms_T_1;
	wire cmd_write_perms = cmd_write | _cmd_write_perms_T_2;
	wire [6:0] _ae_array_T = (misaligned ? eff_array : 7'h00);
	wire [6:0] _ae_array_T_2 = (cmd_lrsc ? 7'h7f : 7'h00);
	wire [6:0] ae_array = _ae_array_T | _ae_array_T_2;
	wire [6:0] _ae_ld_array_T = ~pr_array;
	wire [6:0] _ae_ld_array_T_1 = ae_array | _ae_ld_array_T;
	wire [6:0] ae_ld_array = (cmd_read ? _ae_ld_array_T_1 : 7'h00);
	wire [6:0] _ae_st_array_T = ~pw_array;
	wire [6:0] _ae_st_array_T_1 = ae_array | _ae_st_array_T;
	wire [6:0] _ae_st_array_T_2 = (cmd_write_perms ? _ae_st_array_T_1 : 7'h00);
	wire [6:0] _ae_st_array_T_3 = ~ppp_array;
	wire [6:0] _ae_st_array_T_4 = (cmd_put_partial ? _ae_st_array_T_3 : 7'h00);
	wire [6:0] _ae_st_array_T_5 = _ae_st_array_T_2 | _ae_st_array_T_4;
	wire [6:0] _ae_st_array_T_7 = (cmd_amo_logical ? _ae_st_array_T_3 : 7'h00);
	wire [6:0] _ae_st_array_T_8 = _ae_st_array_T_5 | _ae_st_array_T_7;
	wire [6:0] _ae_st_array_T_10 = (cmd_amo_arithmetic ? _ae_st_array_T_3 : 7'h00);
	wire [6:0] ae_st_array = _ae_st_array_T_8 | _ae_st_array_T_10;
	wire [6:0] pf_ld_array = (cmd_read ? 7'h3f : 7'h00);
	wire [6:0] pf_st_array = (cmd_write_perms ? 7'h3f : 7'h00);
	wire [6:0] _io_resp_pf_ld_T_1 = pf_ld_array & 7'h40;
	wire [6:0] _io_resp_pf_st_T_1 = pf_st_array & 7'h40;
	wire [6:0] _io_resp_ae_ld_T = ae_ld_array & 7'h40;
	wire [6:0] _io_resp_ae_st_T = ae_st_array & 7'h40;
	PMPChecker pmp(
		.io_prv(pmp_io_prv),
		.io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
		.io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
		.io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
		.io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
		.io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
		.io_pmp_0_addr(pmp_io_pmp_0_addr),
		.io_pmp_0_mask(pmp_io_pmp_0_mask),
		.io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
		.io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
		.io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
		.io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
		.io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
		.io_pmp_1_addr(pmp_io_pmp_1_addr),
		.io_pmp_1_mask(pmp_io_pmp_1_mask),
		.io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
		.io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
		.io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
		.io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
		.io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
		.io_pmp_2_addr(pmp_io_pmp_2_addr),
		.io_pmp_2_mask(pmp_io_pmp_2_mask),
		.io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
		.io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
		.io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
		.io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
		.io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
		.io_pmp_3_addr(pmp_io_pmp_3_addr),
		.io_pmp_3_mask(pmp_io_pmp_3_mask),
		.io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
		.io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
		.io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
		.io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
		.io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
		.io_pmp_4_addr(pmp_io_pmp_4_addr),
		.io_pmp_4_mask(pmp_io_pmp_4_mask),
		.io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
		.io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
		.io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
		.io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
		.io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
		.io_pmp_5_addr(pmp_io_pmp_5_addr),
		.io_pmp_5_mask(pmp_io_pmp_5_mask),
		.io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
		.io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
		.io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
		.io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
		.io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
		.io_pmp_6_addr(pmp_io_pmp_6_addr),
		.io_pmp_6_mask(pmp_io_pmp_6_mask),
		.io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
		.io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
		.io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
		.io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
		.io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
		.io_pmp_7_addr(pmp_io_pmp_7_addr),
		.io_pmp_7_mask(pmp_io_pmp_7_mask),
		.io_addr(pmp_io_addr),
		.io_r(pmp_io_r),
		.io_w(pmp_io_w),
		.io_x(pmp_io_x)
	);
	assign io_resp_paddr = {vpn, io_req_bits_vaddr[11:0]};
	assign io_resp_pf_ld = |_io_resp_pf_ld_T_1;
	assign io_resp_pf_st = |_io_resp_pf_st_T_1;
	assign io_resp_ae_ld = |_io_resp_ae_ld_T;
	assign io_resp_ae_st = |_io_resp_ae_st_T;
	assign io_resp_ma_ld = misaligned & cmd_read;
	assign io_resp_ma_st = misaligned & cmd_write;
	assign pmp_io_prv = mpu_priv[1:0];
	assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l;
	assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a;
	assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x;
	assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w;
	assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r;
	assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr;
	assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask;
	assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l;
	assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a;
	assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x;
	assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w;
	assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r;
	assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr;
	assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask;
	assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l;
	assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a;
	assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x;
	assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w;
	assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r;
	assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr;
	assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask;
	assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l;
	assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a;
	assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x;
	assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w;
	assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r;
	assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr;
	assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask;
	assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l;
	assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a;
	assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x;
	assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w;
	assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r;
	assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr;
	assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask;
	assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l;
	assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a;
	assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x;
	assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w;
	assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r;
	assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr;
	assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask;
	assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l;
	assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a;
	assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x;
	assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w;
	assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r;
	assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr;
	assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask;
	assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l;
	assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a;
	assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x;
	assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w;
	assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r;
	assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr;
	assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask;
	assign pmp_io_addr = {mpu_ppn, io_req_bits_vaddr[11:0]};
endmodule
module DCacheModuleImpl_Anon_1 (
	io_in_2_valid,
	io_in_2_bits_addr,
	io_in_3_valid,
	io_in_3_bits_addr,
	io_in_5_ready,
	io_in_5_valid,
	io_in_7_ready,
	io_in_7_valid,
	io_in_7_bits_addr,
	io_out_valid,
	io_out_bits_write,
	io_out_bits_addr
);
	input io_in_2_valid;
	input [31:0] io_in_2_bits_addr;
	input io_in_3_valid;
	input [31:0] io_in_3_bits_addr;
	output wire io_in_5_ready;
	input io_in_5_valid;
	output wire io_in_7_ready;
	input io_in_7_valid;
	input [31:0] io_in_7_bits_addr;
	output wire io_out_valid;
	output wire io_out_bits_write;
	output wire [31:0] io_out_bits_addr;
	wire [31:0] _GEN_22 = (io_in_3_valid ? io_in_3_bits_addr : io_in_7_bits_addr);
	wire _GEN_29 = io_in_2_valid | io_in_3_valid;
	wire grant_4 = ~_GEN_29;
	assign io_in_5_ready = ~_GEN_29;
	assign io_in_7_ready = ~_GEN_29;
	assign io_out_valid = ~grant_4 | io_in_7_valid;
	assign io_out_bits_write = io_in_2_valid | io_in_3_valid;
	assign io_out_bits_addr = (io_in_2_valid ? io_in_2_bits_addr : _GEN_22);
endmodule
module DCacheDataArray (
	clock,
	io_req_valid,
	io_req_bits_addr,
	io_req_bits_write,
	io_req_bits_wdata,
	io_req_bits_eccMask,
	io_resp_0
);
	input clock;
	input io_req_valid;
	input [13:0] io_req_bits_addr;
	input io_req_bits_write;
	input [31:0] io_req_bits_wdata;
	input [3:0] io_req_bits_eccMask;
	output wire [31:0] io_resp_0;
	wire [11:0] data_arrays_0_RW0_addr;
	wire data_arrays_0_RW0_en;
	wire data_arrays_0_RW0_clk;
	wire data_arrays_0_RW0_wmode;
	wire [7:0] data_arrays_0_RW0_wdata_0;
	wire [7:0] data_arrays_0_RW0_wdata_1;
	wire [7:0] data_arrays_0_RW0_wdata_2;
	wire [7:0] data_arrays_0_RW0_wdata_3;
	wire [7:0] data_arrays_0_RW0_rdata_0;
	wire [7:0] data_arrays_0_RW0_rdata_1;
	wire [7:0] data_arrays_0_RW0_rdata_2;
	wire [7:0] data_arrays_0_RW0_rdata_3;
	wire data_arrays_0_RW0_wmask_0;
	wire data_arrays_0_RW0_wmask_1;
	wire data_arrays_0_RW0_wmask_2;
	wire data_arrays_0_RW0_wmask_3;
	wire _rdata_T = io_req_valid & io_req_bits_write;
	wire _rdata_data_T_1 = io_req_valid & ~io_req_bits_write;
	wire [15:0] rdata_lo = {data_arrays_0_RW0_rdata_1, data_arrays_0_RW0_rdata_0};
	wire [15:0] rdata_hi = {data_arrays_0_RW0_rdata_3, data_arrays_0_RW0_rdata_2};
	data_arrays_0 data_arrays_0(
		.RW0_addr(data_arrays_0_RW0_addr),
		.RW0_en(data_arrays_0_RW0_en),
		.RW0_clk(data_arrays_0_RW0_clk),
		.RW0_wmode(data_arrays_0_RW0_wmode),
		.RW0_wdata_0(data_arrays_0_RW0_wdata_0),
		.RW0_wdata_1(data_arrays_0_RW0_wdata_1),
		.RW0_wdata_2(data_arrays_0_RW0_wdata_2),
		.RW0_wdata_3(data_arrays_0_RW0_wdata_3),
		.RW0_rdata_0(data_arrays_0_RW0_rdata_0),
		.RW0_rdata_1(data_arrays_0_RW0_rdata_1),
		.RW0_rdata_2(data_arrays_0_RW0_rdata_2),
		.RW0_rdata_3(data_arrays_0_RW0_rdata_3),
		.RW0_wmask_0(data_arrays_0_RW0_wmask_0),
		.RW0_wmask_1(data_arrays_0_RW0_wmask_1),
		.RW0_wmask_2(data_arrays_0_RW0_wmask_2),
		.RW0_wmask_3(data_arrays_0_RW0_wmask_3)
	);
	assign io_resp_0 = {rdata_hi, rdata_lo};
	assign data_arrays_0_RW0_clk = clock;
	assign data_arrays_0_RW0_wdata_0 = io_req_bits_wdata[7:0];
	assign data_arrays_0_RW0_wdata_1 = io_req_bits_wdata[15:8];
	assign data_arrays_0_RW0_wdata_2 = io_req_bits_wdata[23:16];
	assign data_arrays_0_RW0_wdata_3 = io_req_bits_wdata[31:24];
	assign data_arrays_0_RW0_wmask_0 = io_req_bits_eccMask[0];
	assign data_arrays_0_RW0_wmask_1 = io_req_bits_eccMask[1];
	assign data_arrays_0_RW0_wmask_2 = io_req_bits_eccMask[2];
	assign data_arrays_0_RW0_wmask_3 = io_req_bits_eccMask[3];
	assign data_arrays_0_RW0_en = _rdata_data_T_1 | _rdata_T;
	assign data_arrays_0_RW0_wmode = io_req_bits_write;
	assign data_arrays_0_RW0_addr = io_req_bits_addr[13:2];
endmodule
module DCacheModuleImpl_Anon_2 (
	io_in_0_valid,
	io_in_0_bits_addr,
	io_in_0_bits_write,
	io_in_0_bits_wdata,
	io_in_0_bits_eccMask,
	io_in_1_ready,
	io_in_1_valid,
	io_in_1_bits_addr,
	io_in_1_bits_write,
	io_in_1_bits_wdata,
	io_in_1_bits_eccMask,
	io_in_3_ready,
	io_in_3_valid,
	io_in_3_bits_addr,
	io_in_3_bits_wdata,
	io_in_3_bits_wordMask,
	io_out_valid,
	io_out_bits_addr,
	io_out_bits_write,
	io_out_bits_wdata,
	io_out_bits_eccMask
);
	input io_in_0_valid;
	input [13:0] io_in_0_bits_addr;
	input io_in_0_bits_write;
	input [31:0] io_in_0_bits_wdata;
	input [3:0] io_in_0_bits_eccMask;
	output wire io_in_1_ready;
	input io_in_1_valid;
	input [13:0] io_in_1_bits_addr;
	input io_in_1_bits_write;
	input [31:0] io_in_1_bits_wdata;
	input [3:0] io_in_1_bits_eccMask;
	output wire io_in_3_ready;
	input io_in_3_valid;
	input [13:0] io_in_3_bits_addr;
	input [31:0] io_in_3_bits_wdata;
	input io_in_3_bits_wordMask;
	output wire io_out_valid;
	output wire [13:0] io_out_bits_addr;
	output wire io_out_bits_write;
	output wire [31:0] io_out_bits_wdata;
	output wire [3:0] io_out_bits_eccMask;
	wire [3:0] _GEN_9 = (io_in_1_valid ? io_in_1_bits_eccMask : 4'hf);
	wire [31:0] _GEN_11 = (io_in_1_valid ? io_in_1_bits_wdata : io_in_3_bits_wdata);
	wire [13:0] _GEN_13 = (io_in_1_valid ? io_in_1_bits_addr : io_in_3_bits_addr);
	wire grant_2 = ~(io_in_0_valid | io_in_1_valid);
	assign io_in_1_ready = ~io_in_0_valid;
	assign io_in_3_ready = ~(io_in_0_valid | io_in_1_valid);
	assign io_out_valid = ~grant_2 | io_in_3_valid;
	assign io_out_bits_addr = (io_in_0_valid ? io_in_0_bits_addr : _GEN_13);
	assign io_out_bits_write = (io_in_0_valid ? io_in_0_bits_write : io_in_1_valid & io_in_1_bits_write);
	assign io_out_bits_wdata = (io_in_0_valid ? io_in_0_bits_wdata : _GEN_11);
	assign io_out_bits_eccMask = (io_in_0_valid ? io_in_0_bits_eccMask : _GEN_9);
endmodule
module AMOALU (
	io_cmd,
	io_lhs,
	io_rhs,
	io_out_unmasked
);
	input [4:0] io_cmd;
	input [31:0] io_lhs;
	input [31:0] io_rhs;
	output wire [31:0] io_out_unmasked;
	wire max = (io_cmd == 5'h0d) | (io_cmd == 5'h0f);
	wire min = (io_cmd == 5'h0c) | (io_cmd == 5'h0e);
	wire add = io_cmd == 5'h08;
	wire _logic_and_T = io_cmd == 5'h0a;
	wire logic_and = (io_cmd == 5'h0a) | (io_cmd == 5'h0b);
	wire logic_xor = (io_cmd == 5'h09) | _logic_and_T;
	wire [31:0] adder_out = io_lhs + io_rhs;
	wire [4:0] _less_signed_T = io_cmd & 5'h02;
	wire less_signed = _less_signed_T == 5'h00;
	wire _less_T_6 = io_lhs < io_rhs;
	wire _less_T_9 = (less_signed ? io_lhs[31] : io_rhs[31]);
	wire less = (io_lhs[31] == io_rhs[31] ? _less_T_6 : _less_T_9);
	wire _minmax_T = (less ? min : max);
	wire [31:0] minmax = (_minmax_T ? io_lhs : io_rhs);
	wire [31:0] _logic_T = io_lhs & io_rhs;
	wire [31:0] _logic_T_1 = (logic_and ? _logic_T : 32'h00000000);
	wire [31:0] _logic_T_2 = io_lhs ^ io_rhs;
	wire [31:0] _logic_T_3 = (logic_xor ? _logic_T_2 : 32'h00000000);
	wire [31:0] logic_ = _logic_T_1 | _logic_T_3;
	wire [31:0] _out_T_1 = (logic_and | logic_xor ? logic_ : minmax);
	assign io_out_unmasked = (add ? adder_out : _out_T_1);
endmodule
module DCache (
	clock,
	reset,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	io_cpu_req_ready,
	io_cpu_req_valid,
	io_cpu_req_bits_addr,
	io_cpu_req_bits_tag,
	io_cpu_req_bits_cmd,
	io_cpu_req_bits_size,
	io_cpu_req_bits_signed,
	io_cpu_req_bits_dprv,
	io_cpu_req_bits_no_xcpt,
	io_cpu_s1_kill,
	io_cpu_s1_data_data,
	io_cpu_s1_data_mask,
	io_cpu_s2_nack,
	io_cpu_resp_valid,
	io_cpu_resp_bits_addr,
	io_cpu_resp_bits_tag,
	io_cpu_resp_bits_cmd,
	io_cpu_resp_bits_size,
	io_cpu_resp_bits_signed,
	io_cpu_resp_bits_dprv,
	io_cpu_resp_bits_dv,
	io_cpu_resp_bits_data,
	io_cpu_resp_bits_mask,
	io_cpu_resp_bits_replay,
	io_cpu_resp_bits_has_data,
	io_cpu_resp_bits_data_word_bypass,
	io_cpu_resp_bits_data_raw,
	io_cpu_resp_bits_store_data,
	io_cpu_replay_next,
	io_cpu_s2_xcpt_ma_ld,
	io_cpu_s2_xcpt_ma_st,
	io_cpu_s2_xcpt_pf_ld,
	io_cpu_s2_xcpt_pf_st,
	io_cpu_s2_xcpt_gf_ld,
	io_cpu_s2_xcpt_gf_st,
	io_cpu_s2_xcpt_ae_ld,
	io_cpu_s2_xcpt_ae_st,
	io_cpu_ordered,
	io_cpu_perf_grant,
	io_ptw_status_debug,
	io_ptw_pmp_0_cfg_l,
	io_ptw_pmp_0_cfg_a,
	io_ptw_pmp_0_cfg_x,
	io_ptw_pmp_0_cfg_w,
	io_ptw_pmp_0_cfg_r,
	io_ptw_pmp_0_addr,
	io_ptw_pmp_0_mask,
	io_ptw_pmp_1_cfg_l,
	io_ptw_pmp_1_cfg_a,
	io_ptw_pmp_1_cfg_x,
	io_ptw_pmp_1_cfg_w,
	io_ptw_pmp_1_cfg_r,
	io_ptw_pmp_1_addr,
	io_ptw_pmp_1_mask,
	io_ptw_pmp_2_cfg_l,
	io_ptw_pmp_2_cfg_a,
	io_ptw_pmp_2_cfg_x,
	io_ptw_pmp_2_cfg_w,
	io_ptw_pmp_2_cfg_r,
	io_ptw_pmp_2_addr,
	io_ptw_pmp_2_mask,
	io_ptw_pmp_3_cfg_l,
	io_ptw_pmp_3_cfg_a,
	io_ptw_pmp_3_cfg_x,
	io_ptw_pmp_3_cfg_w,
	io_ptw_pmp_3_cfg_r,
	io_ptw_pmp_3_addr,
	io_ptw_pmp_3_mask,
	io_ptw_pmp_4_cfg_l,
	io_ptw_pmp_4_cfg_a,
	io_ptw_pmp_4_cfg_x,
	io_ptw_pmp_4_cfg_w,
	io_ptw_pmp_4_cfg_r,
	io_ptw_pmp_4_addr,
	io_ptw_pmp_4_mask,
	io_ptw_pmp_5_cfg_l,
	io_ptw_pmp_5_cfg_a,
	io_ptw_pmp_5_cfg_x,
	io_ptw_pmp_5_cfg_w,
	io_ptw_pmp_5_cfg_r,
	io_ptw_pmp_5_addr,
	io_ptw_pmp_5_mask,
	io_ptw_pmp_6_cfg_l,
	io_ptw_pmp_6_cfg_a,
	io_ptw_pmp_6_cfg_x,
	io_ptw_pmp_6_cfg_w,
	io_ptw_pmp_6_cfg_r,
	io_ptw_pmp_6_addr,
	io_ptw_pmp_6_mask,
	io_ptw_pmp_7_cfg_l,
	io_ptw_pmp_7_cfg_a,
	io_ptw_pmp_7_cfg_x,
	io_ptw_pmp_7_cfg_w,
	io_ptw_pmp_7_cfg_r,
	io_ptw_pmp_7_addr,
	io_ptw_pmp_7_mask
);
	input clock;
	input reset;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [3:0] auto_out_d_bits_size;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	output wire io_cpu_req_ready;
	input io_cpu_req_valid;
	input [31:0] io_cpu_req_bits_addr;
	input [6:0] io_cpu_req_bits_tag;
	input [4:0] io_cpu_req_bits_cmd;
	input [1:0] io_cpu_req_bits_size;
	input io_cpu_req_bits_signed;
	input [1:0] io_cpu_req_bits_dprv;
	input io_cpu_req_bits_no_xcpt;
	input io_cpu_s1_kill;
	input [31:0] io_cpu_s1_data_data;
	input [3:0] io_cpu_s1_data_mask;
	output wire io_cpu_s2_nack;
	output wire io_cpu_resp_valid;
	output wire [31:0] io_cpu_resp_bits_addr;
	output wire [6:0] io_cpu_resp_bits_tag;
	output wire [4:0] io_cpu_resp_bits_cmd;
	output wire [1:0] io_cpu_resp_bits_size;
	output wire io_cpu_resp_bits_signed;
	output wire [1:0] io_cpu_resp_bits_dprv;
	output wire io_cpu_resp_bits_dv;
	output wire [31:0] io_cpu_resp_bits_data;
	output wire [3:0] io_cpu_resp_bits_mask;
	output wire io_cpu_resp_bits_replay;
	output wire io_cpu_resp_bits_has_data;
	output wire [31:0] io_cpu_resp_bits_data_word_bypass;
	output wire [31:0] io_cpu_resp_bits_data_raw;
	output wire [31:0] io_cpu_resp_bits_store_data;
	output wire io_cpu_replay_next;
	output wire io_cpu_s2_xcpt_ma_ld;
	output wire io_cpu_s2_xcpt_ma_st;
	output wire io_cpu_s2_xcpt_pf_ld;
	output wire io_cpu_s2_xcpt_pf_st;
	output wire io_cpu_s2_xcpt_gf_ld;
	output wire io_cpu_s2_xcpt_gf_st;
	output wire io_cpu_s2_xcpt_ae_ld;
	output wire io_cpu_s2_xcpt_ae_st;
	output wire io_cpu_ordered;
	output wire io_cpu_perf_grant;
	input io_ptw_status_debug;
	input io_ptw_pmp_0_cfg_l;
	input [1:0] io_ptw_pmp_0_cfg_a;
	input io_ptw_pmp_0_cfg_x;
	input io_ptw_pmp_0_cfg_w;
	input io_ptw_pmp_0_cfg_r;
	input [29:0] io_ptw_pmp_0_addr;
	input [31:0] io_ptw_pmp_0_mask;
	input io_ptw_pmp_1_cfg_l;
	input [1:0] io_ptw_pmp_1_cfg_a;
	input io_ptw_pmp_1_cfg_x;
	input io_ptw_pmp_1_cfg_w;
	input io_ptw_pmp_1_cfg_r;
	input [29:0] io_ptw_pmp_1_addr;
	input [31:0] io_ptw_pmp_1_mask;
	input io_ptw_pmp_2_cfg_l;
	input [1:0] io_ptw_pmp_2_cfg_a;
	input io_ptw_pmp_2_cfg_x;
	input io_ptw_pmp_2_cfg_w;
	input io_ptw_pmp_2_cfg_r;
	input [29:0] io_ptw_pmp_2_addr;
	input [31:0] io_ptw_pmp_2_mask;
	input io_ptw_pmp_3_cfg_l;
	input [1:0] io_ptw_pmp_3_cfg_a;
	input io_ptw_pmp_3_cfg_x;
	input io_ptw_pmp_3_cfg_w;
	input io_ptw_pmp_3_cfg_r;
	input [29:0] io_ptw_pmp_3_addr;
	input [31:0] io_ptw_pmp_3_mask;
	input io_ptw_pmp_4_cfg_l;
	input [1:0] io_ptw_pmp_4_cfg_a;
	input io_ptw_pmp_4_cfg_x;
	input io_ptw_pmp_4_cfg_w;
	input io_ptw_pmp_4_cfg_r;
	input [29:0] io_ptw_pmp_4_addr;
	input [31:0] io_ptw_pmp_4_mask;
	input io_ptw_pmp_5_cfg_l;
	input [1:0] io_ptw_pmp_5_cfg_a;
	input io_ptw_pmp_5_cfg_x;
	input io_ptw_pmp_5_cfg_w;
	input io_ptw_pmp_5_cfg_r;
	input [29:0] io_ptw_pmp_5_addr;
	input [31:0] io_ptw_pmp_5_mask;
	input io_ptw_pmp_6_cfg_l;
	input [1:0] io_ptw_pmp_6_cfg_a;
	input io_ptw_pmp_6_cfg_x;
	input io_ptw_pmp_6_cfg_w;
	input io_ptw_pmp_6_cfg_r;
	input [29:0] io_ptw_pmp_6_addr;
	input [31:0] io_ptw_pmp_6_mask;
	input io_ptw_pmp_7_cfg_l;
	input [1:0] io_ptw_pmp_7_cfg_a;
	input io_ptw_pmp_7_cfg_x;
	input io_ptw_pmp_7_cfg_w;
	input io_ptw_pmp_7_cfg_r;
	input [29:0] io_ptw_pmp_7_addr;
	input [31:0] io_ptw_pmp_7_mask;
	wire tlb_io_req_valid;
	wire [31:0] tlb_io_req_bits_vaddr;
	wire [1:0] tlb_io_req_bits_size;
	wire [4:0] tlb_io_req_bits_cmd;
	wire [1:0] tlb_io_req_bits_prv;
	wire [31:0] tlb_io_resp_paddr;
	wire tlb_io_resp_pf_ld;
	wire tlb_io_resp_pf_st;
	wire tlb_io_resp_ae_ld;
	wire tlb_io_resp_ae_st;
	wire tlb_io_resp_ma_ld;
	wire tlb_io_resp_ma_st;
	wire tlb_io_ptw_status_debug;
	wire tlb_io_ptw_pmp_0_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_0_cfg_a;
	wire tlb_io_ptw_pmp_0_cfg_x;
	wire tlb_io_ptw_pmp_0_cfg_w;
	wire tlb_io_ptw_pmp_0_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_0_addr;
	wire [31:0] tlb_io_ptw_pmp_0_mask;
	wire tlb_io_ptw_pmp_1_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_1_cfg_a;
	wire tlb_io_ptw_pmp_1_cfg_x;
	wire tlb_io_ptw_pmp_1_cfg_w;
	wire tlb_io_ptw_pmp_1_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_1_addr;
	wire [31:0] tlb_io_ptw_pmp_1_mask;
	wire tlb_io_ptw_pmp_2_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_2_cfg_a;
	wire tlb_io_ptw_pmp_2_cfg_x;
	wire tlb_io_ptw_pmp_2_cfg_w;
	wire tlb_io_ptw_pmp_2_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_2_addr;
	wire [31:0] tlb_io_ptw_pmp_2_mask;
	wire tlb_io_ptw_pmp_3_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_3_cfg_a;
	wire tlb_io_ptw_pmp_3_cfg_x;
	wire tlb_io_ptw_pmp_3_cfg_w;
	wire tlb_io_ptw_pmp_3_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_3_addr;
	wire [31:0] tlb_io_ptw_pmp_3_mask;
	wire tlb_io_ptw_pmp_4_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_4_cfg_a;
	wire tlb_io_ptw_pmp_4_cfg_x;
	wire tlb_io_ptw_pmp_4_cfg_w;
	wire tlb_io_ptw_pmp_4_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_4_addr;
	wire [31:0] tlb_io_ptw_pmp_4_mask;
	wire tlb_io_ptw_pmp_5_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_5_cfg_a;
	wire tlb_io_ptw_pmp_5_cfg_x;
	wire tlb_io_ptw_pmp_5_cfg_w;
	wire tlb_io_ptw_pmp_5_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_5_addr;
	wire [31:0] tlb_io_ptw_pmp_5_mask;
	wire tlb_io_ptw_pmp_6_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_6_cfg_a;
	wire tlb_io_ptw_pmp_6_cfg_x;
	wire tlb_io_ptw_pmp_6_cfg_w;
	wire tlb_io_ptw_pmp_6_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_6_addr;
	wire [31:0] tlb_io_ptw_pmp_6_mask;
	wire tlb_io_ptw_pmp_7_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_7_cfg_a;
	wire tlb_io_ptw_pmp_7_cfg_x;
	wire tlb_io_ptw_pmp_7_cfg_w;
	wire tlb_io_ptw_pmp_7_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_7_addr;
	wire [31:0] tlb_io_ptw_pmp_7_mask;
	wire pma_checker_io_req_valid;
	wire [31:0] pma_checker_io_req_bits_vaddr;
	wire [1:0] pma_checker_io_req_bits_size;
	wire [4:0] pma_checker_io_req_bits_cmd;
	wire [1:0] pma_checker_io_req_bits_prv;
	wire [31:0] pma_checker_io_resp_paddr;
	wire pma_checker_io_resp_pf_ld;
	wire pma_checker_io_resp_pf_st;
	wire pma_checker_io_resp_ae_ld;
	wire pma_checker_io_resp_ae_st;
	wire pma_checker_io_resp_ma_ld;
	wire pma_checker_io_resp_ma_st;
	wire pma_checker_io_ptw_status_debug;
	wire pma_checker_io_ptw_pmp_0_cfg_l;
	wire [1:0] pma_checker_io_ptw_pmp_0_cfg_a;
	wire pma_checker_io_ptw_pmp_0_cfg_x;
	wire pma_checker_io_ptw_pmp_0_cfg_w;
	wire pma_checker_io_ptw_pmp_0_cfg_r;
	wire [29:0] pma_checker_io_ptw_pmp_0_addr;
	wire [31:0] pma_checker_io_ptw_pmp_0_mask;
	wire pma_checker_io_ptw_pmp_1_cfg_l;
	wire [1:0] pma_checker_io_ptw_pmp_1_cfg_a;
	wire pma_checker_io_ptw_pmp_1_cfg_x;
	wire pma_checker_io_ptw_pmp_1_cfg_w;
	wire pma_checker_io_ptw_pmp_1_cfg_r;
	wire [29:0] pma_checker_io_ptw_pmp_1_addr;
	wire [31:0] pma_checker_io_ptw_pmp_1_mask;
	wire pma_checker_io_ptw_pmp_2_cfg_l;
	wire [1:0] pma_checker_io_ptw_pmp_2_cfg_a;
	wire pma_checker_io_ptw_pmp_2_cfg_x;
	wire pma_checker_io_ptw_pmp_2_cfg_w;
	wire pma_checker_io_ptw_pmp_2_cfg_r;
	wire [29:0] pma_checker_io_ptw_pmp_2_addr;
	wire [31:0] pma_checker_io_ptw_pmp_2_mask;
	wire pma_checker_io_ptw_pmp_3_cfg_l;
	wire [1:0] pma_checker_io_ptw_pmp_3_cfg_a;
	wire pma_checker_io_ptw_pmp_3_cfg_x;
	wire pma_checker_io_ptw_pmp_3_cfg_w;
	wire pma_checker_io_ptw_pmp_3_cfg_r;
	wire [29:0] pma_checker_io_ptw_pmp_3_addr;
	wire [31:0] pma_checker_io_ptw_pmp_3_mask;
	wire pma_checker_io_ptw_pmp_4_cfg_l;
	wire [1:0] pma_checker_io_ptw_pmp_4_cfg_a;
	wire pma_checker_io_ptw_pmp_4_cfg_x;
	wire pma_checker_io_ptw_pmp_4_cfg_w;
	wire pma_checker_io_ptw_pmp_4_cfg_r;
	wire [29:0] pma_checker_io_ptw_pmp_4_addr;
	wire [31:0] pma_checker_io_ptw_pmp_4_mask;
	wire pma_checker_io_ptw_pmp_5_cfg_l;
	wire [1:0] pma_checker_io_ptw_pmp_5_cfg_a;
	wire pma_checker_io_ptw_pmp_5_cfg_x;
	wire pma_checker_io_ptw_pmp_5_cfg_w;
	wire pma_checker_io_ptw_pmp_5_cfg_r;
	wire [29:0] pma_checker_io_ptw_pmp_5_addr;
	wire [31:0] pma_checker_io_ptw_pmp_5_mask;
	wire pma_checker_io_ptw_pmp_6_cfg_l;
	wire [1:0] pma_checker_io_ptw_pmp_6_cfg_a;
	wire pma_checker_io_ptw_pmp_6_cfg_x;
	wire pma_checker_io_ptw_pmp_6_cfg_w;
	wire pma_checker_io_ptw_pmp_6_cfg_r;
	wire [29:0] pma_checker_io_ptw_pmp_6_addr;
	wire [31:0] pma_checker_io_ptw_pmp_6_mask;
	wire pma_checker_io_ptw_pmp_7_cfg_l;
	wire [1:0] pma_checker_io_ptw_pmp_7_cfg_a;
	wire pma_checker_io_ptw_pmp_7_cfg_x;
	wire pma_checker_io_ptw_pmp_7_cfg_w;
	wire pma_checker_io_ptw_pmp_7_cfg_r;
	wire [29:0] pma_checker_io_ptw_pmp_7_addr;
	wire [31:0] pma_checker_io_ptw_pmp_7_mask;
	wire metaArb_io_in_2_valid;
	wire [31:0] metaArb_io_in_2_bits_addr;
	wire metaArb_io_in_3_valid;
	wire [31:0] metaArb_io_in_3_bits_addr;
	wire metaArb_io_in_5_ready;
	wire metaArb_io_in_5_valid;
	wire metaArb_io_in_7_ready;
	wire metaArb_io_in_7_valid;
	wire [31:0] metaArb_io_in_7_bits_addr;
	wire metaArb_io_out_valid;
	wire metaArb_io_out_bits_write;
	wire [31:0] metaArb_io_out_bits_addr;
	wire data_clock;
	wire data_io_req_valid;
	wire [13:0] data_io_req_bits_addr;
	wire data_io_req_bits_write;
	wire [31:0] data_io_req_bits_wdata;
	wire [3:0] data_io_req_bits_eccMask;
	wire [31:0] data_io_resp_0;
	wire dataArb_io_in_0_valid;
	wire [13:0] dataArb_io_in_0_bits_addr;
	wire dataArb_io_in_0_bits_write;
	wire [31:0] dataArb_io_in_0_bits_wdata;
	wire [3:0] dataArb_io_in_0_bits_eccMask;
	wire dataArb_io_in_1_ready;
	wire dataArb_io_in_1_valid;
	wire [13:0] dataArb_io_in_1_bits_addr;
	wire dataArb_io_in_1_bits_write;
	wire [31:0] dataArb_io_in_1_bits_wdata;
	wire [3:0] dataArb_io_in_1_bits_eccMask;
	wire dataArb_io_in_3_ready;
	wire dataArb_io_in_3_valid;
	wire [13:0] dataArb_io_in_3_bits_addr;
	wire [31:0] dataArb_io_in_3_bits_wdata;
	wire dataArb_io_in_3_bits_wordMask;
	wire dataArb_io_out_valid;
	wire [13:0] dataArb_io_out_bits_addr;
	wire dataArb_io_out_bits_write;
	wire [31:0] dataArb_io_out_bits_wdata;
	wire [3:0] dataArb_io_out_bits_eccMask;
	wire [4:0] amoalu_io_cmd;
	wire [31:0] amoalu_io_lhs;
	wire [31:0] amoalu_io_rhs;
	wire [31:0] amoalu_io_out_unmasked;
	wire s1_valid_x12 = io_cpu_req_ready & io_cpu_req_valid;
	reg s1_valid;
	wire s1_valid_masked = s1_valid & ~io_cpu_s1_kill;
	reg [4:0] s1_req_cmd;
	wire _s1_read_T = s1_req_cmd == 5'h00;
	wire _s1_read_T_1 = s1_req_cmd == 5'h10;
	wire _s1_read_T_2 = s1_req_cmd == 5'h06;
	wire _s1_read_T_3 = s1_req_cmd == 5'h07;
	wire _s1_read_T_6 = ((_s1_read_T | _s1_read_T_1) | _s1_read_T_2) | _s1_read_T_3;
	wire _s1_read_T_7 = s1_req_cmd == 5'h04;
	wire _s1_read_T_8 = s1_req_cmd == 5'h09;
	wire _s1_read_T_9 = s1_req_cmd == 5'h0a;
	wire _s1_read_T_10 = s1_req_cmd == 5'h0b;
	wire _s1_read_T_13 = ((_s1_read_T_7 | _s1_read_T_8) | _s1_read_T_9) | _s1_read_T_10;
	wire _s1_read_T_14 = s1_req_cmd == 5'h08;
	wire _s1_read_T_15 = s1_req_cmd == 5'h0c;
	wire _s1_read_T_16 = s1_req_cmd == 5'h0d;
	wire _s1_read_T_17 = s1_req_cmd == 5'h0e;
	wire _s1_read_T_18 = s1_req_cmd == 5'h0f;
	wire _s1_read_T_22 = (((_s1_read_T_14 | _s1_read_T_15) | _s1_read_T_16) | _s1_read_T_17) | _s1_read_T_18;
	wire _s1_read_T_23 = _s1_read_T_13 | _s1_read_T_22;
	wire s1_read = _s1_read_T_6 | _s1_read_T_23;
	reg s2_valid;
	reg [4:0] s2_req_cmd;
	wire _s2_write_T_1 = s2_req_cmd == 5'h11;
	wire _s2_write_T_3 = s2_req_cmd == 5'h07;
	wire _s2_write_T_5 = s2_req_cmd == 5'h04;
	wire _s2_write_T_6 = s2_req_cmd == 5'h09;
	wire _s2_write_T_7 = s2_req_cmd == 5'h0a;
	wire _s2_write_T_8 = s2_req_cmd == 5'h0b;
	wire _s2_write_T_11 = ((_s2_write_T_5 | _s2_write_T_6) | _s2_write_T_7) | _s2_write_T_8;
	wire _s2_write_T_12 = s2_req_cmd == 5'h08;
	wire _s2_write_T_13 = s2_req_cmd == 5'h0c;
	wire _s2_write_T_14 = s2_req_cmd == 5'h0d;
	wire _s2_write_T_15 = s2_req_cmd == 5'h0e;
	wire _s2_write_T_16 = s2_req_cmd == 5'h0f;
	wire _s2_write_T_20 = (((_s2_write_T_12 | _s2_write_T_13) | _s2_write_T_14) | _s2_write_T_15) | _s2_write_T_16;
	wire _s2_write_T_21 = _s2_write_T_11 | _s2_write_T_20;
	wire s2_write = (((s2_req_cmd == 5'h01) | (s2_req_cmd == 5'h11)) | (s2_req_cmd == 5'h07)) | _s2_write_T_21;
	reg pstore1_held;
	wire pstore1_valid_likely = (s2_valid & s2_write) | pstore1_held;
	reg [31:0] pstore1_addr;
	reg [31:0] s1_req_addr;
	wire [31:0] s1_vaddr = {s1_req_addr[31:14], s1_req_addr[13:0]};
	wire _s1_write_T_1 = s1_req_cmd == 5'h11;
	wire s1_write = (((s1_req_cmd == 5'h01) | (s1_req_cmd == 5'h11)) | _s1_read_T_3) | _s1_read_T_23;
	reg [3:0] pstore1_mask;
	wire _s1_hazard_T_10 = |pstore1_mask[3];
	wire _s1_hazard_T_9 = |pstore1_mask[2];
	wire _s1_hazard_T_8 = |pstore1_mask[1];
	wire _s1_hazard_T_7 = |pstore1_mask[0];
	wire [3:0] _s1_hazard_T_11 = {_s1_hazard_T_10, _s1_hazard_T_9, _s1_hazard_T_8, _s1_hazard_T_7};
	wire [3:0] _s1_hazard_T_16 = {_s1_hazard_T_11[3], _s1_hazard_T_11[2], _s1_hazard_T_11[1], _s1_hazard_T_11[0]};
	reg [1:0] s1_req_size;
	wire s1_mask_xwr_upper = s1_req_addr[0] | (s1_req_size >= 2'h1);
	wire s1_mask_xwr_lower = (s1_req_addr[0] ? 1'h0 : 1'h1);
	wire [1:0] _s1_mask_xwr_T = {s1_mask_xwr_upper, s1_mask_xwr_lower};
	wire [1:0] _s1_mask_xwr_upper_T_5 = (s1_req_addr[1] ? _s1_mask_xwr_T : 2'h0);
	wire [1:0] _s1_mask_xwr_upper_T_7 = (s1_req_size >= 2'h2 ? 2'h3 : 2'h0);
	wire [1:0] s1_mask_xwr_upper_1 = _s1_mask_xwr_upper_T_5 | _s1_mask_xwr_upper_T_7;
	wire [1:0] s1_mask_xwr_lower_1 = (s1_req_addr[1] ? 2'h0 : _s1_mask_xwr_T);
	wire [3:0] s1_mask_xwr = {s1_mask_xwr_upper_1, s1_mask_xwr_lower_1};
	wire _s1_hazard_T_24 = |s1_mask_xwr[3];
	wire _s1_hazard_T_23 = |s1_mask_xwr[2];
	wire _s1_hazard_T_22 = |s1_mask_xwr[1];
	wire _s1_hazard_T_21 = |s1_mask_xwr[0];
	wire [3:0] _s1_hazard_T_25 = {_s1_hazard_T_24, _s1_hazard_T_23, _s1_hazard_T_22, _s1_hazard_T_21};
	wire [3:0] _s1_hazard_T_30 = {_s1_hazard_T_25[3], _s1_hazard_T_25[2], _s1_hazard_T_25[1], _s1_hazard_T_25[0]};
	wire [3:0] _s1_hazard_T_31 = _s1_hazard_T_16 & _s1_hazard_T_30;
	wire [3:0] _s1_hazard_T_33 = pstore1_mask & s1_mask_xwr;
	wire _s1_hazard_T_35 = (s1_write ? |_s1_hazard_T_31 : |_s1_hazard_T_33);
	wire _s1_hazard_T_36 = (pstore1_addr[13:2] == s1_vaddr[13:2]) & _s1_hazard_T_35;
	reg pstore2_valid;
	reg [31:0] pstore2_addr;
	reg [3:0] mask;
	wire _s1_hazard_T_48 = |mask[3];
	wire _s1_hazard_T_47 = |mask[2];
	wire _s1_hazard_T_46 = |mask[1];
	wire _s1_hazard_T_45 = |mask[0];
	wire [3:0] _s1_hazard_T_49 = {_s1_hazard_T_48, _s1_hazard_T_47, _s1_hazard_T_46, _s1_hazard_T_45};
	wire [3:0] _s1_hazard_T_54 = {_s1_hazard_T_49[3], _s1_hazard_T_49[2], _s1_hazard_T_49[1], _s1_hazard_T_49[0]};
	wire [3:0] _s1_hazard_T_69 = _s1_hazard_T_54 & _s1_hazard_T_30;
	wire [3:0] _s1_hazard_T_71 = mask & s1_mask_xwr;
	wire _s1_hazard_T_73 = (s1_write ? |_s1_hazard_T_69 : |_s1_hazard_T_71);
	wire _s1_hazard_T_74 = (pstore2_addr[13:2] == s1_vaddr[13:2]) & _s1_hazard_T_73;
	wire _s1_hazard_T_75 = pstore2_valid & _s1_hazard_T_74;
	wire s1_hazard = (pstore1_valid_likely & _s1_hazard_T_36) | _s1_hazard_T_75;
	wire s1_raw_hazard = s1_read & s1_hazard;
	wire [7:0] _s2_valid_no_xcpt_T = {io_cpu_s2_xcpt_ma_ld, io_cpu_s2_xcpt_ma_st, io_cpu_s2_xcpt_pf_ld, io_cpu_s2_xcpt_pf_st, io_cpu_s2_xcpt_gf_ld, io_cpu_s2_xcpt_gf_st, io_cpu_s2_xcpt_ae_ld, io_cpu_s2_xcpt_ae_st};
	wire s2_valid_no_xcpt = s2_valid & ~(|_s2_valid_no_xcpt_T);
	reg s2_not_nacked_in_s1;
	wire s2_valid_masked = s2_valid_no_xcpt & s2_not_nacked_in_s1;
	wire _c_cat_T_48 = s2_req_cmd == 5'h06;
	wire _c_cat_T_49 = (s2_write | (s2_req_cmd == 5'h03)) | (s2_req_cmd == 5'h06);
	reg [1:0] s2_hit_state_state;
	wire [3:0] _T_35 = {s2_write, _c_cat_T_49, s2_hit_state_state};
	wire _T_93 = 4'h3 == _T_35;
	wire _T_90 = 4'h2 == _T_35;
	wire _T_87 = 4'h1 == _T_35;
	wire _T_84 = 4'h7 == _T_35;
	wire _T_81 = 4'h6 == _T_35;
	wire _T_78 = 4'hf == _T_35;
	wire _T_75 = 4'he == _T_35;
	wire _T_72 = 4'h0 == _T_35;
	wire _T_69 = 4'h5 == _T_35;
	wire _T_66 = 4'h4 == _T_35;
	wire _T_63 = 4'hd == _T_35;
	wire _T_60 = 4'hc == _T_35;
	wire s2_hit = _T_93 | (_T_90 | (_T_87 | (_T_84 | (_T_81 | (_T_78 | _T_75)))));
	wire s2_valid_hit_maybe_flush_pre_data_ecc_and_waw = s2_valid_masked & s2_hit;
	wire _s2_read_T = s2_req_cmd == 5'h00;
	wire _s2_read_T_1 = s2_req_cmd == 5'h10;
	wire _s2_read_T_6 = ((_s2_read_T | _s2_read_T_1) | _c_cat_T_48) | _s2_write_T_3;
	wire s2_read = _s2_read_T_6 | _s2_write_T_21;
	wire s2_readwrite = s2_read | s2_write;
	wire s2_valid_hit_pre_data_ecc_and_waw = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_readwrite;
	wire [1:0] _T_62 = (_T_60 ? 2'h1 : 2'h0);
	wire [1:0] _T_65 = (_T_63 ? 2'h2 : _T_62);
	wire [1:0] _T_68 = (_T_66 ? 2'h1 : _T_65);
	wire [1:0] _T_71 = (_T_69 ? 2'h2 : _T_68);
	wire [1:0] _T_74 = (_T_72 ? 2'h0 : _T_71);
	wire [1:0] _T_77 = (_T_75 ? 2'h3 : _T_74);
	wire [1:0] _T_80 = (_T_78 ? 2'h3 : _T_77);
	wire [1:0] _T_83 = (_T_81 ? 2'h2 : _T_80);
	wire [1:0] _T_86 = (_T_84 ? 2'h3 : _T_83);
	wire [1:0] _T_89 = (_T_87 ? 2'h1 : _T_86);
	wire [1:0] _T_92 = (_T_90 ? 2'h2 : _T_89);
	wire [1:0] s2_grow_param = (_T_93 ? 2'h3 : _T_92);
	wire _s2_update_meta_T = s2_hit_state_state == s2_grow_param;
	wire s2_update_meta = ~_s2_update_meta_T;
	wire _T_223 = io_cpu_s2_nack | (s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta);
	reg s1_req_no_xcpt;
	wire s1_readwrite = s1_read | s1_write;
	wire s1_flush_line = (s1_req_cmd == 5'h05) & s1_req_size[0];
	wire s1_cmd_uses_tlb = (s1_readwrite | s1_flush_line) | (s1_req_cmd == 5'h17);
	wire s1_nack = (s1_valid & s1_raw_hazard) | _T_223;
	wire _s1_valid_not_nacked_T = ~s1_nack;
	wire s1_valid_not_nacked = s1_valid & ~s1_nack;
	wire s0_clk_en = metaArb_io_out_valid & ~metaArb_io_out_bits_write;
	wire [31:0] s0_req_addr = {metaArb_io_out_bits_addr[31:6], io_cpu_req_bits_addr[5:0]};
	wire _T = ~metaArb_io_in_7_ready;
	reg [6:0] s1_req_tag;
	reg s1_req_signed;
	reg [1:0] s1_req_dprv;
	reg [31:0] s1_tlb_req_vaddr;
	reg [1:0] s1_tlb_req_size;
	reg [4:0] s1_tlb_req_cmd;
	reg [1:0] s1_tlb_req_prv;
	wire s1_sfence = ((s1_req_cmd == 5'h14) | (s1_req_cmd == 5'h15)) | (s1_req_cmd == 5'h16);
	reg s1_flush_valid;
	reg uncachedInFlight_0;
	reg [31:0] uncachedReqs_0_addr;
	reg [6:0] uncachedReqs_0_tag;
	reg [1:0] uncachedReqs_0_size;
	reg uncachedReqs_0_signed;
	wire _s0_read_T = io_cpu_req_bits_cmd == 5'h00;
	wire _s0_read_T_1 = io_cpu_req_bits_cmd == 5'h10;
	wire _s0_read_T_2 = io_cpu_req_bits_cmd == 5'h06;
	wire _s0_read_T_3 = io_cpu_req_bits_cmd == 5'h07;
	wire _s0_read_T_6 = ((_s0_read_T | _s0_read_T_1) | _s0_read_T_2) | _s0_read_T_3;
	wire _s0_read_T_7 = io_cpu_req_bits_cmd == 5'h04;
	wire _s0_read_T_8 = io_cpu_req_bits_cmd == 5'h09;
	wire _s0_read_T_9 = io_cpu_req_bits_cmd == 5'h0a;
	wire _s0_read_T_10 = io_cpu_req_bits_cmd == 5'h0b;
	wire _s0_read_T_13 = ((_s0_read_T_7 | _s0_read_T_8) | _s0_read_T_9) | _s0_read_T_10;
	wire _s0_read_T_14 = io_cpu_req_bits_cmd == 5'h08;
	wire _s0_read_T_15 = io_cpu_req_bits_cmd == 5'h0c;
	wire _s0_read_T_16 = io_cpu_req_bits_cmd == 5'h0d;
	wire _s0_read_T_17 = io_cpu_req_bits_cmd == 5'h0e;
	wire _s0_read_T_18 = io_cpu_req_bits_cmd == 5'h0f;
	wire _s0_read_T_22 = (((_s0_read_T_14 | _s0_read_T_15) | _s0_read_T_16) | _s0_read_T_17) | _s0_read_T_18;
	wire _s0_read_T_23 = _s0_read_T_13 | _s0_read_T_22;
	wire s0_read = _s0_read_T_6 | _s0_read_T_23;
	wire _dataArb_io_in_3_valid_res_T = io_cpu_req_bits_cmd == 5'h01;
	wire _dataArb_io_in_3_valid_res_T_1 = io_cpu_req_bits_cmd == 5'h03;
	wire _dataArb_io_in_3_valid_res_T_2 = _dataArb_io_in_3_valid_res_T | _dataArb_io_in_3_valid_res_T_1;
	wire res = ~_dataArb_io_in_3_valid_res_T_2;
	wire _dataArb_io_in_3_valid_T_26 = io_cpu_req_bits_cmd == 5'h11;
	wire _dataArb_io_in_3_valid_T_47 = ((_dataArb_io_in_3_valid_res_T | (io_cpu_req_bits_cmd == 5'h11)) | _s0_read_T_3) | _s0_read_T_23;
	wire _dataArb_io_in_3_valid_T_51 = _dataArb_io_in_3_valid_T_47 & _dataArb_io_in_3_valid_T_26;
	wire _dataArb_io_in_3_valid_T_52 = s0_read | _dataArb_io_in_3_valid_T_51;
	wire _dataArb_io_in_3_valid_T_56 = ~reset;
	wire _dataArb_io_in_3_valid_T_58 = io_cpu_req_valid & res;
	wire [31:0] _dataArb_io_in_3_bits_addr_T_2 = {io_cpu_req_bits_addr[31:14], io_cpu_req_bits_addr[13:0]};
	wire _GEN_33 = (~dataArb_io_in_3_ready & s0_read ? 1'h0 : _s1_valid_not_nacked_T);
	wire _s1_did_read_T_54 = dataArb_io_in_3_ready & (io_cpu_req_valid & _dataArb_io_in_3_valid_T_52);
	reg s1_did_read;
	reg s1_read_mask;
	wire _GEN_36 = (_T ? 1'h0 : _GEN_33);
	wire [31:0] s1_paddr = {tlb_io_resp_paddr[31:12], s1_req_addr[11:0]};
	wire inScratchpad = (s1_paddr >= 32'h80000000) & (s1_paddr < 32'h80004000);
	wire [31:0] _tl_d_data_encoded_T_4 = {auto_out_d_bits_data[31:24], auto_out_d_bits_data[23:16], auto_out_d_bits_data[15:8], auto_out_d_bits_data[7:0]};
	wire [3:0] _T_27 = ~io_cpu_s1_data_mask;
	wire [3:0] _T_28 = s1_mask_xwr | _T_27;
	wire s2_valid_x44 = s1_valid_masked & ~s1_sfence;
	reg [31:0] s2_req_addr;
	reg [6:0] s2_req_tag;
	reg [1:0] s2_req_size;
	reg s2_req_signed;
	reg [1:0] s2_req_dprv;
	reg s2_req_no_xcpt;
	reg s2_tlb_xcpt_pf_ld;
	reg s2_tlb_xcpt_pf_st;
	reg s2_tlb_xcpt_ae_ld;
	reg s2_tlb_xcpt_ae_st;
	reg s2_tlb_xcpt_ma_ld;
	reg s2_tlb_xcpt_ma_st;
	reg [31:0] s2_uncached_resp_addr;
	wire _T_34 = s1_valid_not_nacked | s1_flush_valid;
	wire [31:0] _GEN_40 = (s1_valid_not_nacked | s1_flush_valid ? s1_paddr : s2_req_addr);
	wire [6:0] _GEN_41 = (s1_valid_not_nacked | s1_flush_valid ? s1_req_tag : s2_req_tag);
	wire [4:0] _GEN_42 = (s1_valid_not_nacked | s1_flush_valid ? s1_req_cmd : s2_req_cmd);
	wire [1:0] _GEN_43 = (s1_valid_not_nacked | s1_flush_valid ? s1_req_size : s2_req_size);
	wire _GEN_44 = (s1_valid_not_nacked | s1_flush_valid ? s1_req_signed : s2_req_signed);
	reg [31:0] s2_vaddr_r;
	wire [31:0] s2_vaddr = {s2_vaddr_r[31:14], s2_req_addr[13:0]};
	reg s2_flush_valid_pre_tag_ecc;
	wire en = s1_valid | io_cpu_replay_next;
	wire word_en = s1_did_read & s1_read_mask;
	wire [31:0] s1_all_data_ways_0 = data_io_resp_0;
	wire s1_word_en = (~io_cpu_replay_next ? word_en : 1'h1);
	wire [1:0] opc = auto_out_d_bits_opcode[1:0];
	wire [1:0] _T_257 = opc & 2'h1;
	wire data_1 = _T_257 == 2'h1;
	reg blockUncachedGrant;
	wire [2:0] _GEN_244 = {1'd0, opc};
	wire grantIsRefill = _GEN_244 == 3'h5;
	wire _T_284 = ~dataArb_io_in_1_ready;
	wire _grantIsCached_T = _GEN_244 == 3'h4;
	wire grantIsCached = _grantIsCached_T | grantIsRefill;
	reg [9:0] counter;
	wire d_first = counter == 10'h000;
	wire _bundleOut_0_d_ready_T_3 = (grantIsCached ? ~d_first : 1'h1);
	wire _GEN_223 = (grantIsRefill & ~dataArb_io_in_1_ready ? 1'h0 : _bundleOut_0_d_ready_T_3);
	wire tl_out__d_ready = (data_1 & (blockUncachedGrant | s1_valid) ? 1'h0 : _GEN_223);
	wire _T_261 = tl_out__d_ready & auto_out_d_valid;
	wire [1:0] _GEN_180 = (data_1 ? 2'h2 : 2'h1);
	wire [1:0] _GEN_202 = (grantIsCached ? 2'h1 : _GEN_180);
	wire [1:0] s1_data_way = (_T_261 ? _GEN_202 : 2'h1);
	wire [1:0] _s2_data_T_1 = (s1_word_en ? s1_data_way : 2'h0);
	wire [31:0] _s2_data_T_4 = (_s2_data_T_1[0] ? s1_all_data_ways_0 : 32'h00000000);
	wire [31:0] _s2_data_T_5 = (_s2_data_T_1[1] ? _tl_d_data_encoded_T_4 : 32'h00000000);
	wire [31:0] _s2_data_T_6 = _s2_data_T_4 | _s2_data_T_5;
	reg [31:0] s2_data;
	wire s2_hit_valid = s2_hit_state_state > 2'h0;
	wire [15:0] s2_data_corrected_lo = {s2_data[15:8], s2_data[7:0]};
	wire [15:0] s2_data_corrected_hi = {s2_data[31:24], s2_data[23:16]};
	wire [31:0] s2_data_corrected = {s2_data[31:24], s2_data[23:16], s2_data[15:8], s2_data[7:0]};
	wire s2_valid_miss = (s2_valid_masked & s2_readwrite) & ~s2_hit;
	wire _s2_valid_cached_miss_T_2 = |uncachedInFlight_0;
	wire s2_valid_cached_miss = 1'h0;
	wire _s2_cannot_victimize_T = ~s2_flush_valid_pre_tag_ecc;
	wire s2_valid_uncached_pending = s2_valid_miss & ~(&uncachedInFlight_0);
	wire [1:0] s2_victim_state_state = (s2_hit_valid ? s2_hit_state_state : 2'h0);
	wire [3:0] _T_163 = {2'h2, s2_victim_state_state};
	wire _T_188 = 4'hb == _T_163;
	wire _T_192 = 4'h4 == _T_163;
	wire _T_193 = (_T_192 ? 1'h0 : _T_188);
	wire _T_196 = 4'h5 == _T_163;
	wire _T_197 = (_T_196 ? 1'h0 : _T_193);
	wire _T_200 = 4'h6 == _T_163;
	wire _T_201 = (_T_200 ? 1'h0 : _T_197);
	wire _T_204 = 4'h7 == _T_163;
	wire _T_208 = 4'h0 == _T_163;
	wire _T_209 = (_T_208 ? 1'h0 : _T_204 | _T_201);
	wire _T_212 = 4'h1 == _T_163;
	wire _T_213 = (_T_212 ? 1'h0 : _T_209);
	wire _T_216 = 4'h2 == _T_163;
	wire _T_217 = (_T_216 ? 1'h0 : _T_213);
	wire _T_220 = 4'h3 == _T_163;
	wire s2_victim_dirty = _T_220 | _T_217;
	wire s2_dont_nack_uncached = s2_valid_uncached_pending & auto_out_a_ready;
	wire _s2_dont_nack_misc_T_10 = s2_req_cmd == 5'h17;
	wire s2_dont_nack_misc = s2_valid_masked & _s2_dont_nack_misc_T_10;
	wire _io_cpu_s2_nack_T_4 = ~s2_valid_hit_pre_data_ecc_and_waw;
	wire _pstore1_cmd_T = s1_valid_not_nacked & s1_write;
	reg [4:0] pstore1_cmd;
	reg [31:0] pstore1_data;
	wire _pstore1_rmw_T_51 = s1_write & _s1_write_T_1;
	wire _pstore1_rmw_T_52 = s1_read | _pstore1_rmw_T_51;
	reg pstore1_rmw_r;
	wire _pstore1_merge_T = s2_valid_hit_pre_data_ecc_and_waw & s2_write;
	wire pstore_drain_opportunistic = ~_dataArb_io_in_3_valid_T_58;
	reg pstore_drain_on_miss_REG;
	wire pstore1_valid = _pstore1_merge_T | pstore1_held;
	wire pstore_drain_structural = (pstore1_valid_likely & pstore2_valid) & ((s1_valid & s1_write) | pstore1_rmw_r);
	wire _pstore_drain_T_10 = ((pstore1_valid & ~pstore1_rmw_r) | pstore2_valid) & (pstore_drain_opportunistic | pstore_drain_on_miss_REG);
	wire pstore_drain = pstore_drain_structural | _pstore_drain_T_10;
	wire _pstore1_held_T_9 = ~pstore_drain;
	wire advance_pstore1 = pstore1_valid & (pstore2_valid == pstore_drain);
	wire [7:0] _pstore1_storegen_data_mask_T_12 = (pstore1_mask[3] ? 8'hff : 8'h00);
	wire [7:0] _pstore1_storegen_data_mask_T_10 = (pstore1_mask[2] ? 8'hff : 8'h00);
	wire [7:0] _pstore1_storegen_data_mask_T_8 = (pstore1_mask[1] ? 8'hff : 8'h00);
	wire [7:0] _pstore1_storegen_data_mask_T_6 = (pstore1_mask[0] ? 8'hff : 8'h00);
	wire [31:0] mask_1 = {_pstore1_storegen_data_mask_T_12, _pstore1_storegen_data_mask_T_10, _pstore1_storegen_data_mask_T_8, _pstore1_storegen_data_mask_T_6};
	wire [31:0] _pstore1_storegen_data_T = amoalu_io_out_unmasked & mask_1;
	wire [31:0] _pstore1_storegen_data_T_1 = ~mask_1;
	wire [31:0] _pstore1_storegen_data_T_2 = s2_data_corrected & _pstore1_storegen_data_T_1;
	wire [31:0] pstore1_storegen_data = _pstore1_storegen_data_T | _pstore1_storegen_data_T_2;
	reg [7:0] pstore2_storegen_data_r;
	reg [7:0] pstore2_storegen_data_r_1;
	reg [7:0] pstore2_storegen_data_r_2;
	reg [7:0] pstore2_storegen_data_r_3;
	wire [31:0] pstore2_storegen_data = {pstore2_storegen_data_r_3, pstore2_storegen_data_r_2, pstore2_storegen_data_r_1, pstore2_storegen_data_r};
	wire [3:0] _pstore2_storegen_mask_mask_T = ~pstore1_mask;
	wire [3:0] _pstore2_storegen_mask_mask_T_2 = ~_pstore2_storegen_mask_mask_T;
	wire [31:0] _dataArb_io_in_0_bits_addr_T = (pstore2_valid ? pstore2_addr : pstore1_addr);
	wire [31:0] _dataArb_io_in_0_bits_wdata_T = (pstore2_valid ? pstore2_storegen_data : pstore1_data);
	wire [15:0] dataArb_io_in_0_bits_wdata_lo = {_dataArb_io_in_0_bits_wdata_T[15:8], _dataArb_io_in_0_bits_wdata_T[7:0]};
	wire [15:0] dataArb_io_in_0_bits_wdata_hi = {_dataArb_io_in_0_bits_wdata_T[31:24], _dataArb_io_in_0_bits_wdata_T[23:16]};
	wire [3:0] _dataArb_io_in_0_bits_eccMask_T = (pstore2_valid ? mask : pstore1_mask);
	wire _dataArb_io_in_0_bits_eccMask_T_5 = |_dataArb_io_in_0_bits_eccMask_T[0];
	wire _dataArb_io_in_0_bits_eccMask_T_6 = |_dataArb_io_in_0_bits_eccMask_T[1];
	wire _dataArb_io_in_0_bits_eccMask_T_7 = |_dataArb_io_in_0_bits_eccMask_T[2];
	wire _dataArb_io_in_0_bits_eccMask_T_8 = |_dataArb_io_in_0_bits_eccMask_T[3];
	wire [1:0] dataArb_io_in_0_bits_eccMask_lo = {_dataArb_io_in_0_bits_eccMask_T_6, _dataArb_io_in_0_bits_eccMask_T_5};
	wire [1:0] dataArb_io_in_0_bits_eccMask_hi = {_dataArb_io_in_0_bits_eccMask_T_8, _dataArb_io_in_0_bits_eccMask_T_7};
	wire _a_source_T = ~uncachedInFlight_0;
	wire [18:0] a_mask = {15'd0, pstore1_mask};
	wire [1:0] _get_a_mask_sizeOH_T_1 = 2'h1 << s2_req_size[0];
	wire [1:0] get_a_mask_sizeOH = _get_a_mask_sizeOH_T_1 | 2'h1;
	wire _get_a_mask_T = s2_req_size >= 2'h2;
	wire get_a_mask_size = get_a_mask_sizeOH[1];
	wire get_a_mask_bit = s2_req_addr[1];
	wire get_a_mask_nbit = ~get_a_mask_bit;
	wire get_a_mask_acc = _get_a_mask_T | (get_a_mask_size & get_a_mask_nbit);
	wire get_a_mask_acc_1 = _get_a_mask_T | (get_a_mask_size & get_a_mask_bit);
	wire get_a_mask_size_1 = get_a_mask_sizeOH[0];
	wire get_a_mask_bit_1 = s2_req_addr[0];
	wire get_a_mask_nbit_1 = ~get_a_mask_bit_1;
	wire get_a_mask_eq_2 = get_a_mask_nbit & get_a_mask_nbit_1;
	wire get_a_mask_acc_2 = get_a_mask_acc | (get_a_mask_size_1 & get_a_mask_eq_2);
	wire get_a_mask_eq_3 = get_a_mask_nbit & get_a_mask_bit_1;
	wire get_a_mask_acc_3 = get_a_mask_acc | (get_a_mask_size_1 & get_a_mask_eq_3);
	wire get_a_mask_eq_4 = get_a_mask_bit & get_a_mask_nbit_1;
	wire get_a_mask_acc_4 = get_a_mask_acc_1 | (get_a_mask_size_1 & get_a_mask_eq_4);
	wire get_a_mask_eq_5 = get_a_mask_bit & get_a_mask_bit_1;
	wire get_a_mask_acc_5 = get_a_mask_acc_1 | (get_a_mask_size_1 & get_a_mask_eq_5);
	wire [3:0] get_mask = {get_a_mask_acc_5, get_a_mask_acc_4, get_a_mask_acc_3, get_a_mask_acc_2};
	wire [2:0] _atomics_T_1_opcode = (5'h04 == s2_req_cmd ? 3'h3 : 3'h0);
	wire [3:0] atomics_a_size = {2'd0, s2_req_size};
	wire [3:0] _atomics_T_1_size = (5'h04 == s2_req_cmd ? atomics_a_size : 4'h0);
	wire [31:0] _atomics_T_1_address = (5'h04 == s2_req_cmd ? s2_req_addr : 32'h00000000);
	wire [3:0] _atomics_T_1_mask = (5'h04 == s2_req_cmd ? get_mask : 4'h0);
	wire [31:0] _atomics_T_1_data = (5'h04 == s2_req_cmd ? pstore1_data : 32'h00000000);
	wire [2:0] _atomics_T_3_opcode = (5'h09 == s2_req_cmd ? 3'h3 : _atomics_T_1_opcode);
	wire [2:0] _atomics_T_3_param = (5'h09 == s2_req_cmd ? 3'h0 : _atomics_T_1_opcode);
	wire [3:0] _atomics_T_3_size = (5'h09 == s2_req_cmd ? atomics_a_size : _atomics_T_1_size);
	wire [31:0] _atomics_T_3_address = (5'h09 == s2_req_cmd ? s2_req_addr : _atomics_T_1_address);
	wire [3:0] _atomics_T_3_mask = (5'h09 == s2_req_cmd ? get_mask : _atomics_T_1_mask);
	wire [31:0] _atomics_T_3_data = (5'h09 == s2_req_cmd ? pstore1_data : _atomics_T_1_data);
	wire [2:0] _atomics_T_5_opcode = (5'h0a == s2_req_cmd ? 3'h3 : _atomics_T_3_opcode);
	wire [2:0] _atomics_T_5_param = (5'h0a == s2_req_cmd ? 3'h1 : _atomics_T_3_param);
	wire [3:0] _atomics_T_5_size = (5'h0a == s2_req_cmd ? atomics_a_size : _atomics_T_3_size);
	wire [31:0] _atomics_T_5_address = (5'h0a == s2_req_cmd ? s2_req_addr : _atomics_T_3_address);
	wire [3:0] _atomics_T_5_mask = (5'h0a == s2_req_cmd ? get_mask : _atomics_T_3_mask);
	wire [31:0] _atomics_T_5_data = (5'h0a == s2_req_cmd ? pstore1_data : _atomics_T_3_data);
	wire [2:0] _atomics_T_7_opcode = (5'h0b == s2_req_cmd ? 3'h3 : _atomics_T_5_opcode);
	wire [2:0] _atomics_T_7_param = (5'h0b == s2_req_cmd ? 3'h2 : _atomics_T_5_param);
	wire [3:0] _atomics_T_7_size = (5'h0b == s2_req_cmd ? atomics_a_size : _atomics_T_5_size);
	wire [31:0] _atomics_T_7_address = (5'h0b == s2_req_cmd ? s2_req_addr : _atomics_T_5_address);
	wire [3:0] _atomics_T_7_mask = (5'h0b == s2_req_cmd ? get_mask : _atomics_T_5_mask);
	wire [31:0] _atomics_T_7_data = (5'h0b == s2_req_cmd ? pstore1_data : _atomics_T_5_data);
	wire [2:0] _atomics_T_9_opcode = (5'h08 == s2_req_cmd ? 3'h2 : _atomics_T_7_opcode);
	wire [2:0] _atomics_T_9_param = (5'h08 == s2_req_cmd ? 3'h4 : _atomics_T_7_param);
	wire [3:0] _atomics_T_9_size = (5'h08 == s2_req_cmd ? atomics_a_size : _atomics_T_7_size);
	wire [31:0] _atomics_T_9_address = (5'h08 == s2_req_cmd ? s2_req_addr : _atomics_T_7_address);
	wire [3:0] _atomics_T_9_mask = (5'h08 == s2_req_cmd ? get_mask : _atomics_T_7_mask);
	wire [31:0] _atomics_T_9_data = (5'h08 == s2_req_cmd ? pstore1_data : _atomics_T_7_data);
	wire [2:0] _atomics_T_11_opcode = (5'h0c == s2_req_cmd ? 3'h2 : _atomics_T_9_opcode);
	wire [2:0] _atomics_T_11_param = (5'h0c == s2_req_cmd ? 3'h0 : _atomics_T_9_param);
	wire [3:0] _atomics_T_11_size = (5'h0c == s2_req_cmd ? atomics_a_size : _atomics_T_9_size);
	wire [31:0] _atomics_T_11_address = (5'h0c == s2_req_cmd ? s2_req_addr : _atomics_T_9_address);
	wire [3:0] _atomics_T_11_mask = (5'h0c == s2_req_cmd ? get_mask : _atomics_T_9_mask);
	wire [31:0] _atomics_T_11_data = (5'h0c == s2_req_cmd ? pstore1_data : _atomics_T_9_data);
	wire [2:0] _atomics_T_13_opcode = (5'h0d == s2_req_cmd ? 3'h2 : _atomics_T_11_opcode);
	wire [2:0] _atomics_T_13_param = (5'h0d == s2_req_cmd ? 3'h1 : _atomics_T_11_param);
	wire [3:0] _atomics_T_13_size = (5'h0d == s2_req_cmd ? atomics_a_size : _atomics_T_11_size);
	wire [31:0] _atomics_T_13_address = (5'h0d == s2_req_cmd ? s2_req_addr : _atomics_T_11_address);
	wire [3:0] _atomics_T_13_mask = (5'h0d == s2_req_cmd ? get_mask : _atomics_T_11_mask);
	wire [31:0] _atomics_T_13_data = (5'h0d == s2_req_cmd ? pstore1_data : _atomics_T_11_data);
	wire [2:0] _atomics_T_15_opcode = (5'h0e == s2_req_cmd ? 3'h2 : _atomics_T_13_opcode);
	wire [2:0] _atomics_T_15_param = (5'h0e == s2_req_cmd ? 3'h2 : _atomics_T_13_param);
	wire [3:0] _atomics_T_15_size = (5'h0e == s2_req_cmd ? atomics_a_size : _atomics_T_13_size);
	wire [31:0] _atomics_T_15_address = (5'h0e == s2_req_cmd ? s2_req_addr : _atomics_T_13_address);
	wire [3:0] _atomics_T_15_mask = (5'h0e == s2_req_cmd ? get_mask : _atomics_T_13_mask);
	wire [31:0] _atomics_T_15_data = (5'h0e == s2_req_cmd ? pstore1_data : _atomics_T_13_data);
	wire [2:0] atomics_opcode = (5'h0f == s2_req_cmd ? 3'h2 : _atomics_T_15_opcode);
	wire [2:0] atomics_param = (5'h0f == s2_req_cmd ? 3'h3 : _atomics_T_15_param);
	wire [3:0] atomics_size = (5'h0f == s2_req_cmd ? atomics_a_size : _atomics_T_15_size);
	wire [31:0] atomics_address = (5'h0f == s2_req_cmd ? s2_req_addr : _atomics_T_15_address);
	wire [3:0] atomics_mask = (5'h0f == s2_req_cmd ? get_mask : _atomics_T_15_mask);
	wire [31:0] atomics_data = (5'h0f == s2_req_cmd ? pstore1_data : _atomics_T_15_data);
	wire _tl_out_a_valid_T_10 = ~s2_victim_dirty;
	wire _tl_out_a_valid_T_12 = 1'h0 & _tl_out_a_valid_T_10;
	wire tl_out_a_valid = s2_valid_uncached_pending | _tl_out_a_valid_T_12;
	wire [2:0] _tl_out_a_bits_T_4_opcode = (~s2_read ? 3'h0 : atomics_opcode);
	wire [2:0] _tl_out_a_bits_T_4_param = (~s2_read ? 3'h0 : atomics_param);
	wire [3:0] _tl_out_a_bits_T_4_size = (~s2_read ? atomics_a_size : atomics_size);
	wire [31:0] _tl_out_a_bits_T_4_address = (~s2_read ? s2_req_addr : atomics_address);
	wire [3:0] _tl_out_a_bits_T_4_mask = (~s2_read ? get_mask : atomics_mask);
	wire [31:0] _tl_out_a_bits_T_4_data = (~s2_read ? pstore1_data : atomics_data);
	wire [2:0] _tl_out_a_bits_T_5_opcode = (_s2_write_T_1 ? 3'h1 : _tl_out_a_bits_T_4_opcode);
	wire [2:0] _tl_out_a_bits_T_5_param = (_s2_write_T_1 ? 3'h0 : _tl_out_a_bits_T_4_param);
	wire [3:0] _tl_out_a_bits_T_5_size = (_s2_write_T_1 ? atomics_a_size : _tl_out_a_bits_T_4_size);
	wire [31:0] _tl_out_a_bits_T_5_address = (_s2_write_T_1 ? s2_req_addr : _tl_out_a_bits_T_4_address);
	wire [3:0] putpartial_mask = a_mask[3:0];
	wire [3:0] _tl_out_a_bits_T_5_mask = (_s2_write_T_1 ? putpartial_mask : _tl_out_a_bits_T_4_mask);
	wire [31:0] _tl_out_a_bits_T_5_data = (_s2_write_T_1 ? pstore1_data : _tl_out_a_bits_T_4_data);
	wire _T_244 = auto_out_a_ready & tl_out_a_valid;
	wire _GEN_158 = _T_244 | uncachedInFlight_0;
	wire [26:0] _beats1_decode_T_1 = 27'h0000fff << auto_out_d_bits_size;
	wire [11:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[11:0];
	wire [9:0] beats1_decode = _beats1_decode_T_3[11:2];
	wire beats1_opdata = auto_out_d_bits_opcode[0];
	wire [9:0] beats1 = (beats1_opdata ? beats1_decode : 10'h000);
	wire [9:0] counter1 = counter - 10'h001;
	wire d_last = (counter == 10'h001) | (beats1 == 10'h000);
	wire d_done = d_last & _T_261;
	wire _T_248 = auto_out_d_bits_opcode == 3'h1;
	wire _T_249 = auto_out_d_bits_opcode == 3'h0;
	wire _T_250 = auto_out_d_bits_opcode == 3'h2;
	wire _T_252 = (_T_248 | _T_249) | _T_250;
	wire [31:0] dontCareBits = {s1_paddr[31:2], 2'h0};
	wire [31:0] _GEN_249 = {30'd0, uncachedReqs_0_addr[1:0]};
	wire [31:0] _s2_req_addr_T_1 = dontCareBits | _GEN_249;
	wire _GEN_224 = (auto_out_d_valid ? 1'h0 : _GEN_36);
	wire _GEN_225 = auto_out_d_valid | (auto_out_d_valid & grantIsRefill);
	wire _GEN_226 = (auto_out_d_valid ? 1'h0 : dataArb_io_in_0_bits_write);
	wire _io_cpu_ordered_T = ~s1_req_no_xcpt;
	reg io_cpu_s2_xcpt_REG;
	wire _T_299 = _c_cat_T_48 | _s2_write_T_3;
	reg doUncachedResp;
	wire [15:0] io_cpu_resp_bits_data_shifted = (get_a_mask_bit ? s2_data_corrected[31:16] : s2_data_corrected[15:0]);
	wire _io_cpu_resp_bits_data_T_3 = s2_req_signed & io_cpu_resp_bits_data_shifted[15];
	wire [15:0] _io_cpu_resp_bits_data_T_5 = (_io_cpu_resp_bits_data_T_3 ? 16'hffff : 16'h0000);
	wire [15:0] _io_cpu_resp_bits_data_T_7 = (s2_req_size == 2'h1 ? _io_cpu_resp_bits_data_T_5 : s2_data_corrected[31:16]);
	wire [31:0] _io_cpu_resp_bits_data_T_8 = {_io_cpu_resp_bits_data_T_7, io_cpu_resp_bits_data_shifted};
	wire [7:0] io_cpu_resp_bits_data_shifted_1 = (get_a_mask_bit_1 ? _io_cpu_resp_bits_data_T_8[15:8] : _io_cpu_resp_bits_data_T_8[7:0]);
	wire _io_cpu_resp_bits_data_T_12 = s2_req_signed & io_cpu_resp_bits_data_shifted_1[7];
	wire [23:0] _io_cpu_resp_bits_data_T_14 = (_io_cpu_resp_bits_data_T_12 ? 24'hffffff : 24'h000000);
	wire [23:0] _io_cpu_resp_bits_data_T_16 = (s2_req_size == 2'h0 ? _io_cpu_resp_bits_data_T_14 : _io_cpu_resp_bits_data_T_8[31:8]);
	wire _s1_flush_valid_T = metaArb_io_in_5_ready & metaArb_io_in_5_valid;
	wire _T_314 = ~grantIsCached;
	TLB tlb(
		.io_req_valid(tlb_io_req_valid),
		.io_req_bits_vaddr(tlb_io_req_bits_vaddr),
		.io_req_bits_size(tlb_io_req_bits_size),
		.io_req_bits_cmd(tlb_io_req_bits_cmd),
		.io_req_bits_prv(tlb_io_req_bits_prv),
		.io_resp_paddr(tlb_io_resp_paddr),
		.io_resp_pf_ld(tlb_io_resp_pf_ld),
		.io_resp_pf_st(tlb_io_resp_pf_st),
		.io_resp_ae_ld(tlb_io_resp_ae_ld),
		.io_resp_ae_st(tlb_io_resp_ae_st),
		.io_resp_ma_ld(tlb_io_resp_ma_ld),
		.io_resp_ma_st(tlb_io_resp_ma_st),
		.io_ptw_status_debug(tlb_io_ptw_status_debug),
		.io_ptw_pmp_0_cfg_l(tlb_io_ptw_pmp_0_cfg_l),
		.io_ptw_pmp_0_cfg_a(tlb_io_ptw_pmp_0_cfg_a),
		.io_ptw_pmp_0_cfg_x(tlb_io_ptw_pmp_0_cfg_x),
		.io_ptw_pmp_0_cfg_w(tlb_io_ptw_pmp_0_cfg_w),
		.io_ptw_pmp_0_cfg_r(tlb_io_ptw_pmp_0_cfg_r),
		.io_ptw_pmp_0_addr(tlb_io_ptw_pmp_0_addr),
		.io_ptw_pmp_0_mask(tlb_io_ptw_pmp_0_mask),
		.io_ptw_pmp_1_cfg_l(tlb_io_ptw_pmp_1_cfg_l),
		.io_ptw_pmp_1_cfg_a(tlb_io_ptw_pmp_1_cfg_a),
		.io_ptw_pmp_1_cfg_x(tlb_io_ptw_pmp_1_cfg_x),
		.io_ptw_pmp_1_cfg_w(tlb_io_ptw_pmp_1_cfg_w),
		.io_ptw_pmp_1_cfg_r(tlb_io_ptw_pmp_1_cfg_r),
		.io_ptw_pmp_1_addr(tlb_io_ptw_pmp_1_addr),
		.io_ptw_pmp_1_mask(tlb_io_ptw_pmp_1_mask),
		.io_ptw_pmp_2_cfg_l(tlb_io_ptw_pmp_2_cfg_l),
		.io_ptw_pmp_2_cfg_a(tlb_io_ptw_pmp_2_cfg_a),
		.io_ptw_pmp_2_cfg_x(tlb_io_ptw_pmp_2_cfg_x),
		.io_ptw_pmp_2_cfg_w(tlb_io_ptw_pmp_2_cfg_w),
		.io_ptw_pmp_2_cfg_r(tlb_io_ptw_pmp_2_cfg_r),
		.io_ptw_pmp_2_addr(tlb_io_ptw_pmp_2_addr),
		.io_ptw_pmp_2_mask(tlb_io_ptw_pmp_2_mask),
		.io_ptw_pmp_3_cfg_l(tlb_io_ptw_pmp_3_cfg_l),
		.io_ptw_pmp_3_cfg_a(tlb_io_ptw_pmp_3_cfg_a),
		.io_ptw_pmp_3_cfg_x(tlb_io_ptw_pmp_3_cfg_x),
		.io_ptw_pmp_3_cfg_w(tlb_io_ptw_pmp_3_cfg_w),
		.io_ptw_pmp_3_cfg_r(tlb_io_ptw_pmp_3_cfg_r),
		.io_ptw_pmp_3_addr(tlb_io_ptw_pmp_3_addr),
		.io_ptw_pmp_3_mask(tlb_io_ptw_pmp_3_mask),
		.io_ptw_pmp_4_cfg_l(tlb_io_ptw_pmp_4_cfg_l),
		.io_ptw_pmp_4_cfg_a(tlb_io_ptw_pmp_4_cfg_a),
		.io_ptw_pmp_4_cfg_x(tlb_io_ptw_pmp_4_cfg_x),
		.io_ptw_pmp_4_cfg_w(tlb_io_ptw_pmp_4_cfg_w),
		.io_ptw_pmp_4_cfg_r(tlb_io_ptw_pmp_4_cfg_r),
		.io_ptw_pmp_4_addr(tlb_io_ptw_pmp_4_addr),
		.io_ptw_pmp_4_mask(tlb_io_ptw_pmp_4_mask),
		.io_ptw_pmp_5_cfg_l(tlb_io_ptw_pmp_5_cfg_l),
		.io_ptw_pmp_5_cfg_a(tlb_io_ptw_pmp_5_cfg_a),
		.io_ptw_pmp_5_cfg_x(tlb_io_ptw_pmp_5_cfg_x),
		.io_ptw_pmp_5_cfg_w(tlb_io_ptw_pmp_5_cfg_w),
		.io_ptw_pmp_5_cfg_r(tlb_io_ptw_pmp_5_cfg_r),
		.io_ptw_pmp_5_addr(tlb_io_ptw_pmp_5_addr),
		.io_ptw_pmp_5_mask(tlb_io_ptw_pmp_5_mask),
		.io_ptw_pmp_6_cfg_l(tlb_io_ptw_pmp_6_cfg_l),
		.io_ptw_pmp_6_cfg_a(tlb_io_ptw_pmp_6_cfg_a),
		.io_ptw_pmp_6_cfg_x(tlb_io_ptw_pmp_6_cfg_x),
		.io_ptw_pmp_6_cfg_w(tlb_io_ptw_pmp_6_cfg_w),
		.io_ptw_pmp_6_cfg_r(tlb_io_ptw_pmp_6_cfg_r),
		.io_ptw_pmp_6_addr(tlb_io_ptw_pmp_6_addr),
		.io_ptw_pmp_6_mask(tlb_io_ptw_pmp_6_mask),
		.io_ptw_pmp_7_cfg_l(tlb_io_ptw_pmp_7_cfg_l),
		.io_ptw_pmp_7_cfg_a(tlb_io_ptw_pmp_7_cfg_a),
		.io_ptw_pmp_7_cfg_x(tlb_io_ptw_pmp_7_cfg_x),
		.io_ptw_pmp_7_cfg_w(tlb_io_ptw_pmp_7_cfg_w),
		.io_ptw_pmp_7_cfg_r(tlb_io_ptw_pmp_7_cfg_r),
		.io_ptw_pmp_7_addr(tlb_io_ptw_pmp_7_addr),
		.io_ptw_pmp_7_mask(tlb_io_ptw_pmp_7_mask)
	);
	TLB pma_checker(
		.io_req_valid(pma_checker_io_req_valid),
		.io_req_bits_vaddr(pma_checker_io_req_bits_vaddr),
		.io_req_bits_size(pma_checker_io_req_bits_size),
		.io_req_bits_cmd(pma_checker_io_req_bits_cmd),
		.io_req_bits_prv(pma_checker_io_req_bits_prv),
		.io_resp_paddr(pma_checker_io_resp_paddr),
		.io_resp_pf_ld(pma_checker_io_resp_pf_ld),
		.io_resp_pf_st(pma_checker_io_resp_pf_st),
		.io_resp_ae_ld(pma_checker_io_resp_ae_ld),
		.io_resp_ae_st(pma_checker_io_resp_ae_st),
		.io_resp_ma_ld(pma_checker_io_resp_ma_ld),
		.io_resp_ma_st(pma_checker_io_resp_ma_st),
		.io_ptw_status_debug(pma_checker_io_ptw_status_debug),
		.io_ptw_pmp_0_cfg_l(pma_checker_io_ptw_pmp_0_cfg_l),
		.io_ptw_pmp_0_cfg_a(pma_checker_io_ptw_pmp_0_cfg_a),
		.io_ptw_pmp_0_cfg_x(pma_checker_io_ptw_pmp_0_cfg_x),
		.io_ptw_pmp_0_cfg_w(pma_checker_io_ptw_pmp_0_cfg_w),
		.io_ptw_pmp_0_cfg_r(pma_checker_io_ptw_pmp_0_cfg_r),
		.io_ptw_pmp_0_addr(pma_checker_io_ptw_pmp_0_addr),
		.io_ptw_pmp_0_mask(pma_checker_io_ptw_pmp_0_mask),
		.io_ptw_pmp_1_cfg_l(pma_checker_io_ptw_pmp_1_cfg_l),
		.io_ptw_pmp_1_cfg_a(pma_checker_io_ptw_pmp_1_cfg_a),
		.io_ptw_pmp_1_cfg_x(pma_checker_io_ptw_pmp_1_cfg_x),
		.io_ptw_pmp_1_cfg_w(pma_checker_io_ptw_pmp_1_cfg_w),
		.io_ptw_pmp_1_cfg_r(pma_checker_io_ptw_pmp_1_cfg_r),
		.io_ptw_pmp_1_addr(pma_checker_io_ptw_pmp_1_addr),
		.io_ptw_pmp_1_mask(pma_checker_io_ptw_pmp_1_mask),
		.io_ptw_pmp_2_cfg_l(pma_checker_io_ptw_pmp_2_cfg_l),
		.io_ptw_pmp_2_cfg_a(pma_checker_io_ptw_pmp_2_cfg_a),
		.io_ptw_pmp_2_cfg_x(pma_checker_io_ptw_pmp_2_cfg_x),
		.io_ptw_pmp_2_cfg_w(pma_checker_io_ptw_pmp_2_cfg_w),
		.io_ptw_pmp_2_cfg_r(pma_checker_io_ptw_pmp_2_cfg_r),
		.io_ptw_pmp_2_addr(pma_checker_io_ptw_pmp_2_addr),
		.io_ptw_pmp_2_mask(pma_checker_io_ptw_pmp_2_mask),
		.io_ptw_pmp_3_cfg_l(pma_checker_io_ptw_pmp_3_cfg_l),
		.io_ptw_pmp_3_cfg_a(pma_checker_io_ptw_pmp_3_cfg_a),
		.io_ptw_pmp_3_cfg_x(pma_checker_io_ptw_pmp_3_cfg_x),
		.io_ptw_pmp_3_cfg_w(pma_checker_io_ptw_pmp_3_cfg_w),
		.io_ptw_pmp_3_cfg_r(pma_checker_io_ptw_pmp_3_cfg_r),
		.io_ptw_pmp_3_addr(pma_checker_io_ptw_pmp_3_addr),
		.io_ptw_pmp_3_mask(pma_checker_io_ptw_pmp_3_mask),
		.io_ptw_pmp_4_cfg_l(pma_checker_io_ptw_pmp_4_cfg_l),
		.io_ptw_pmp_4_cfg_a(pma_checker_io_ptw_pmp_4_cfg_a),
		.io_ptw_pmp_4_cfg_x(pma_checker_io_ptw_pmp_4_cfg_x),
		.io_ptw_pmp_4_cfg_w(pma_checker_io_ptw_pmp_4_cfg_w),
		.io_ptw_pmp_4_cfg_r(pma_checker_io_ptw_pmp_4_cfg_r),
		.io_ptw_pmp_4_addr(pma_checker_io_ptw_pmp_4_addr),
		.io_ptw_pmp_4_mask(pma_checker_io_ptw_pmp_4_mask),
		.io_ptw_pmp_5_cfg_l(pma_checker_io_ptw_pmp_5_cfg_l),
		.io_ptw_pmp_5_cfg_a(pma_checker_io_ptw_pmp_5_cfg_a),
		.io_ptw_pmp_5_cfg_x(pma_checker_io_ptw_pmp_5_cfg_x),
		.io_ptw_pmp_5_cfg_w(pma_checker_io_ptw_pmp_5_cfg_w),
		.io_ptw_pmp_5_cfg_r(pma_checker_io_ptw_pmp_5_cfg_r),
		.io_ptw_pmp_5_addr(pma_checker_io_ptw_pmp_5_addr),
		.io_ptw_pmp_5_mask(pma_checker_io_ptw_pmp_5_mask),
		.io_ptw_pmp_6_cfg_l(pma_checker_io_ptw_pmp_6_cfg_l),
		.io_ptw_pmp_6_cfg_a(pma_checker_io_ptw_pmp_6_cfg_a),
		.io_ptw_pmp_6_cfg_x(pma_checker_io_ptw_pmp_6_cfg_x),
		.io_ptw_pmp_6_cfg_w(pma_checker_io_ptw_pmp_6_cfg_w),
		.io_ptw_pmp_6_cfg_r(pma_checker_io_ptw_pmp_6_cfg_r),
		.io_ptw_pmp_6_addr(pma_checker_io_ptw_pmp_6_addr),
		.io_ptw_pmp_6_mask(pma_checker_io_ptw_pmp_6_mask),
		.io_ptw_pmp_7_cfg_l(pma_checker_io_ptw_pmp_7_cfg_l),
		.io_ptw_pmp_7_cfg_a(pma_checker_io_ptw_pmp_7_cfg_a),
		.io_ptw_pmp_7_cfg_x(pma_checker_io_ptw_pmp_7_cfg_x),
		.io_ptw_pmp_7_cfg_w(pma_checker_io_ptw_pmp_7_cfg_w),
		.io_ptw_pmp_7_cfg_r(pma_checker_io_ptw_pmp_7_cfg_r),
		.io_ptw_pmp_7_addr(pma_checker_io_ptw_pmp_7_addr),
		.io_ptw_pmp_7_mask(pma_checker_io_ptw_pmp_7_mask)
	);
	DCacheModuleImpl_Anon_1 metaArb(
		.io_in_2_valid(metaArb_io_in_2_valid),
		.io_in_2_bits_addr(metaArb_io_in_2_bits_addr),
		.io_in_3_valid(metaArb_io_in_3_valid),
		.io_in_3_bits_addr(metaArb_io_in_3_bits_addr),
		.io_in_5_ready(metaArb_io_in_5_ready),
		.io_in_5_valid(metaArb_io_in_5_valid),
		.io_in_7_ready(metaArb_io_in_7_ready),
		.io_in_7_valid(metaArb_io_in_7_valid),
		.io_in_7_bits_addr(metaArb_io_in_7_bits_addr),
		.io_out_valid(metaArb_io_out_valid),
		.io_out_bits_write(metaArb_io_out_bits_write),
		.io_out_bits_addr(metaArb_io_out_bits_addr)
	);
	DCacheDataArray data(
		.clock(data_clock),
		.io_req_valid(data_io_req_valid),
		.io_req_bits_addr(data_io_req_bits_addr),
		.io_req_bits_write(data_io_req_bits_write),
		.io_req_bits_wdata(data_io_req_bits_wdata),
		.io_req_bits_eccMask(data_io_req_bits_eccMask),
		.io_resp_0(data_io_resp_0)
	);
	DCacheModuleImpl_Anon_2 dataArb(
		.io_in_0_valid(dataArb_io_in_0_valid),
		.io_in_0_bits_addr(dataArb_io_in_0_bits_addr),
		.io_in_0_bits_write(dataArb_io_in_0_bits_write),
		.io_in_0_bits_wdata(dataArb_io_in_0_bits_wdata),
		.io_in_0_bits_eccMask(dataArb_io_in_0_bits_eccMask),
		.io_in_1_ready(dataArb_io_in_1_ready),
		.io_in_1_valid(dataArb_io_in_1_valid),
		.io_in_1_bits_addr(dataArb_io_in_1_bits_addr),
		.io_in_1_bits_write(dataArb_io_in_1_bits_write),
		.io_in_1_bits_wdata(dataArb_io_in_1_bits_wdata),
		.io_in_1_bits_eccMask(dataArb_io_in_1_bits_eccMask),
		.io_in_3_ready(dataArb_io_in_3_ready),
		.io_in_3_valid(dataArb_io_in_3_valid),
		.io_in_3_bits_addr(dataArb_io_in_3_bits_addr),
		.io_in_3_bits_wdata(dataArb_io_in_3_bits_wdata),
		.io_in_3_bits_wordMask(dataArb_io_in_3_bits_wordMask),
		.io_out_valid(dataArb_io_out_valid),
		.io_out_bits_addr(dataArb_io_out_bits_addr),
		.io_out_bits_write(dataArb_io_out_bits_write),
		.io_out_bits_wdata(dataArb_io_out_bits_wdata),
		.io_out_bits_eccMask(dataArb_io_out_bits_eccMask)
	);
	AMOALU amoalu(
		.io_cmd(amoalu_io_cmd),
		.io_lhs(amoalu_io_lhs),
		.io_rhs(amoalu_io_rhs),
		.io_out_unmasked(amoalu_io_out_unmasked)
	);
	assign auto_out_a_valid = s2_valid_uncached_pending | _tl_out_a_valid_T_12;
	assign auto_out_a_bits_opcode = (~s2_write ? 3'h4 : _tl_out_a_bits_T_5_opcode);
	assign auto_out_a_bits_param = (~s2_write ? 3'h0 : _tl_out_a_bits_T_5_param);
	assign auto_out_a_bits_size = (~s2_write ? atomics_a_size : _tl_out_a_bits_T_5_size);
	assign auto_out_a_bits_address = (~s2_write ? s2_req_addr : _tl_out_a_bits_T_5_address);
	assign auto_out_a_bits_mask = (~s2_write ? get_mask : _tl_out_a_bits_T_5_mask);
	assign auto_out_a_bits_data = (~s2_write ? 32'h00000000 : _tl_out_a_bits_T_5_data);
	assign auto_out_d_ready = (data_1 & (blockUncachedGrant | s1_valid) ? 1'h0 : _GEN_223);
	assign io_cpu_req_ready = (data_1 & (blockUncachedGrant | s1_valid) ? _GEN_224 : _GEN_36);
	assign io_cpu_s2_nack = ((s2_valid_no_xcpt & ~s2_dont_nack_uncached) & ~s2_dont_nack_misc) & ~s2_valid_hit_pre_data_ecc_and_waw;
	assign io_cpu_resp_valid = s2_valid_hit_pre_data_ecc_and_waw | doUncachedResp;
	assign io_cpu_resp_bits_addr = (doUncachedResp ? s2_uncached_resp_addr : s2_req_addr);
	assign io_cpu_resp_bits_tag = s2_req_tag;
	assign io_cpu_resp_bits_cmd = s2_req_cmd;
	assign io_cpu_resp_bits_size = s2_req_size;
	assign io_cpu_resp_bits_signed = s2_req_signed;
	assign io_cpu_resp_bits_dprv = s2_req_dprv;
	assign io_cpu_resp_bits_dv = 1'h0;
	assign io_cpu_resp_bits_data = {_io_cpu_resp_bits_data_T_16, io_cpu_resp_bits_data_shifted_1};
	assign io_cpu_resp_bits_mask = 4'h0;
	assign io_cpu_resp_bits_replay = doUncachedResp;
	assign io_cpu_resp_bits_has_data = _s2_read_T_6 | _s2_write_T_21;
	assign io_cpu_resp_bits_data_word_bypass = {s2_data_corrected_hi, s2_data_corrected_lo};
	assign io_cpu_resp_bits_data_raw = {s2_data_corrected_hi, s2_data_corrected_lo};
	assign io_cpu_resp_bits_store_data = pstore1_data;
	assign io_cpu_replay_next = _T_261 & data_1;
	assign io_cpu_s2_xcpt_ma_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ma_ld;
	assign io_cpu_s2_xcpt_ma_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ma_st;
	assign io_cpu_s2_xcpt_pf_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_pf_ld;
	assign io_cpu_s2_xcpt_pf_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_pf_st;
	assign io_cpu_s2_xcpt_gf_ld = 1'h0;
	assign io_cpu_s2_xcpt_gf_st = 1'h0;
	assign io_cpu_s2_xcpt_ae_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ae_ld;
	assign io_cpu_s2_xcpt_ae_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ae_st;
	assign io_cpu_ordered = ~(((s1_valid & ~s1_req_no_xcpt) | (s2_valid & ~s2_req_no_xcpt)) | _s2_valid_cached_miss_T_2);
	assign io_cpu_perf_grant = auto_out_d_valid & d_last;
	assign tlb_io_req_valid = s1_valid_masked & s1_cmd_uses_tlb;
	assign tlb_io_req_bits_vaddr = s1_tlb_req_vaddr;
	assign tlb_io_req_bits_size = s1_tlb_req_size;
	assign tlb_io_req_bits_cmd = s1_tlb_req_cmd;
	assign tlb_io_req_bits_prv = s1_tlb_req_prv;
	assign tlb_io_ptw_status_debug = io_ptw_status_debug;
	assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l;
	assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a;
	assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x;
	assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w;
	assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r;
	assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr;
	assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask;
	assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l;
	assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a;
	assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x;
	assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w;
	assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r;
	assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr;
	assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask;
	assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l;
	assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a;
	assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x;
	assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w;
	assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r;
	assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr;
	assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask;
	assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l;
	assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a;
	assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x;
	assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w;
	assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r;
	assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr;
	assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask;
	assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l;
	assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a;
	assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x;
	assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w;
	assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r;
	assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr;
	assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask;
	assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l;
	assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a;
	assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x;
	assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w;
	assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r;
	assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr;
	assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask;
	assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l;
	assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a;
	assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x;
	assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w;
	assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r;
	assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr;
	assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask;
	assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l;
	assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a;
	assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x;
	assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w;
	assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r;
	assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr;
	assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask;
	assign pma_checker_io_req_valid = 1'h0;
	assign pma_checker_io_req_bits_vaddr = 32'h00000000;
	assign pma_checker_io_req_bits_size = s1_req_size;
	assign pma_checker_io_req_bits_cmd = s1_req_cmd;
	assign pma_checker_io_req_bits_prv = 2'h0;
	assign pma_checker_io_ptw_status_debug = 1'h0;
	assign pma_checker_io_ptw_pmp_0_cfg_l = 1'h0;
	assign pma_checker_io_ptw_pmp_0_cfg_a = 2'h0;
	assign pma_checker_io_ptw_pmp_0_cfg_x = 1'h0;
	assign pma_checker_io_ptw_pmp_0_cfg_w = 1'h0;
	assign pma_checker_io_ptw_pmp_0_cfg_r = 1'h0;
	assign pma_checker_io_ptw_pmp_0_addr = 30'h00000000;
	assign pma_checker_io_ptw_pmp_0_mask = 32'h00000000;
	assign pma_checker_io_ptw_pmp_1_cfg_l = 1'h0;
	assign pma_checker_io_ptw_pmp_1_cfg_a = 2'h0;
	assign pma_checker_io_ptw_pmp_1_cfg_x = 1'h0;
	assign pma_checker_io_ptw_pmp_1_cfg_w = 1'h0;
	assign pma_checker_io_ptw_pmp_1_cfg_r = 1'h0;
	assign pma_checker_io_ptw_pmp_1_addr = 30'h00000000;
	assign pma_checker_io_ptw_pmp_1_mask = 32'h00000000;
	assign pma_checker_io_ptw_pmp_2_cfg_l = 1'h0;
	assign pma_checker_io_ptw_pmp_2_cfg_a = 2'h0;
	assign pma_checker_io_ptw_pmp_2_cfg_x = 1'h0;
	assign pma_checker_io_ptw_pmp_2_cfg_w = 1'h0;
	assign pma_checker_io_ptw_pmp_2_cfg_r = 1'h0;
	assign pma_checker_io_ptw_pmp_2_addr = 30'h00000000;
	assign pma_checker_io_ptw_pmp_2_mask = 32'h00000000;
	assign pma_checker_io_ptw_pmp_3_cfg_l = 1'h0;
	assign pma_checker_io_ptw_pmp_3_cfg_a = 2'h0;
	assign pma_checker_io_ptw_pmp_3_cfg_x = 1'h0;
	assign pma_checker_io_ptw_pmp_3_cfg_w = 1'h0;
	assign pma_checker_io_ptw_pmp_3_cfg_r = 1'h0;
	assign pma_checker_io_ptw_pmp_3_addr = 30'h00000000;
	assign pma_checker_io_ptw_pmp_3_mask = 32'h00000000;
	assign pma_checker_io_ptw_pmp_4_cfg_l = 1'h0;
	assign pma_checker_io_ptw_pmp_4_cfg_a = 2'h0;
	assign pma_checker_io_ptw_pmp_4_cfg_x = 1'h0;
	assign pma_checker_io_ptw_pmp_4_cfg_w = 1'h0;
	assign pma_checker_io_ptw_pmp_4_cfg_r = 1'h0;
	assign pma_checker_io_ptw_pmp_4_addr = 30'h00000000;
	assign pma_checker_io_ptw_pmp_4_mask = 32'h00000000;
	assign pma_checker_io_ptw_pmp_5_cfg_l = 1'h0;
	assign pma_checker_io_ptw_pmp_5_cfg_a = 2'h0;
	assign pma_checker_io_ptw_pmp_5_cfg_x = 1'h0;
	assign pma_checker_io_ptw_pmp_5_cfg_w = 1'h0;
	assign pma_checker_io_ptw_pmp_5_cfg_r = 1'h0;
	assign pma_checker_io_ptw_pmp_5_addr = 30'h00000000;
	assign pma_checker_io_ptw_pmp_5_mask = 32'h00000000;
	assign pma_checker_io_ptw_pmp_6_cfg_l = 1'h0;
	assign pma_checker_io_ptw_pmp_6_cfg_a = 2'h0;
	assign pma_checker_io_ptw_pmp_6_cfg_x = 1'h0;
	assign pma_checker_io_ptw_pmp_6_cfg_w = 1'h0;
	assign pma_checker_io_ptw_pmp_6_cfg_r = 1'h0;
	assign pma_checker_io_ptw_pmp_6_addr = 30'h00000000;
	assign pma_checker_io_ptw_pmp_6_mask = 32'h00000000;
	assign pma_checker_io_ptw_pmp_7_cfg_l = 1'h0;
	assign pma_checker_io_ptw_pmp_7_cfg_a = 2'h0;
	assign pma_checker_io_ptw_pmp_7_cfg_x = 1'h0;
	assign pma_checker_io_ptw_pmp_7_cfg_w = 1'h0;
	assign pma_checker_io_ptw_pmp_7_cfg_r = 1'h0;
	assign pma_checker_io_ptw_pmp_7_addr = 30'h00000000;
	assign pma_checker_io_ptw_pmp_7_mask = 32'h00000000;
	assign metaArb_io_in_2_valid = s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta;
	assign metaArb_io_in_2_bits_addr = {io_cpu_req_bits_addr[31:14], s2_vaddr[13:0]};
	assign metaArb_io_in_3_valid = (grantIsCached & d_done) & ~auto_out_d_bits_denied;
	assign metaArb_io_in_3_bits_addr = {io_cpu_req_bits_addr[31:14], s2_vaddr[13:0]};
	assign metaArb_io_in_5_valid = 1'h0;
	assign metaArb_io_in_7_valid = io_cpu_req_valid;
	assign metaArb_io_in_7_bits_addr = io_cpu_req_bits_addr;
	assign data_clock = clock;
	assign data_io_req_valid = dataArb_io_out_valid;
	assign data_io_req_bits_addr = dataArb_io_out_bits_addr;
	assign data_io_req_bits_write = dataArb_io_out_bits_write;
	assign data_io_req_bits_wdata = dataArb_io_out_bits_wdata;
	assign data_io_req_bits_eccMask = dataArb_io_out_bits_eccMask;
	assign dataArb_io_in_0_valid = pstore_drain_structural | _pstore_drain_T_10;
	assign dataArb_io_in_0_bits_addr = _dataArb_io_in_0_bits_addr_T[13:0];
	assign dataArb_io_in_0_bits_write = pstore_drain_structural | _pstore_drain_T_10;
	assign dataArb_io_in_0_bits_wdata = {dataArb_io_in_0_bits_wdata_hi, dataArb_io_in_0_bits_wdata_lo};
	assign dataArb_io_in_0_bits_eccMask = {dataArb_io_in_0_bits_eccMask_hi, dataArb_io_in_0_bits_eccMask_lo};
	assign dataArb_io_in_1_valid = (data_1 & (blockUncachedGrant | s1_valid) ? _GEN_225 : auto_out_d_valid & grantIsRefill);
	assign dataArb_io_in_1_bits_addr = dataArb_io_in_0_bits_addr;
	assign dataArb_io_in_1_bits_write = (data_1 & (blockUncachedGrant | s1_valid) ? _GEN_226 : dataArb_io_in_0_bits_write);
	assign dataArb_io_in_1_bits_wdata = dataArb_io_in_0_bits_wdata;
	assign dataArb_io_in_1_bits_eccMask = dataArb_io_in_0_bits_eccMask;
	assign dataArb_io_in_3_valid = io_cpu_req_valid & res;
	assign dataArb_io_in_3_bits_addr = _dataArb_io_in_3_bits_addr_T_2[13:0];
	assign dataArb_io_in_3_bits_wdata = dataArb_io_in_1_bits_wdata;
	assign dataArb_io_in_3_bits_wordMask = 1'h1;
	assign amoalu_io_cmd = pstore1_cmd;
	assign amoalu_io_lhs = {s2_data_corrected_hi, s2_data_corrected_lo};
	assign amoalu_io_rhs = pstore1_data;
	always @(posedge clock) begin
		if (reset)
			s1_valid <= 1'h0;
		else
			s1_valid <= s1_valid_x12;
		if (s0_clk_en)
			s1_req_cmd <= io_cpu_req_bits_cmd;
		if (reset)
			s2_valid <= 1'h0;
		else
			s2_valid <= s2_valid_x44;
		if (_T_261) begin
			if (grantIsCached)
				s2_req_cmd <= _GEN_42;
			else if (data_1)
				s2_req_cmd <= 5'h00;
			else
				s2_req_cmd <= _GEN_42;
		end
		else
			s2_req_cmd <= _GEN_42;
		if (reset)
			pstore1_held <= 1'h0;
		else
			pstore1_held <= (pstore1_valid & pstore2_valid) & ~pstore_drain;
		if (_pstore1_cmd_T)
			pstore1_addr <= s1_vaddr;
		if (s0_clk_en)
			s1_req_addr <= s0_req_addr;
		if (_pstore1_cmd_T)
			if (_s1_write_T_1)
				pstore1_mask <= io_cpu_s1_data_mask;
			else
				pstore1_mask <= s1_mask_xwr;
		if (s0_clk_en)
			s1_req_size <= io_cpu_req_bits_size;
		if (reset)
			pstore2_valid <= 1'h0;
		else
			pstore2_valid <= (pstore2_valid & _pstore1_held_T_9) | advance_pstore1;
		if (advance_pstore1)
			pstore2_addr <= pstore1_addr;
		if (advance_pstore1)
			mask <= _pstore2_storegen_mask_mask_T_2;
		s2_not_nacked_in_s1 <= ~s1_nack;
		if (_T_34)
			if (inScratchpad)
				s2_hit_state_state <= 2'h3;
			else
				s2_hit_state_state <= 2'h0;
		if (s0_clk_en)
			s1_req_no_xcpt <= io_cpu_req_bits_no_xcpt;
		if (s0_clk_en)
			s1_req_tag <= io_cpu_req_bits_tag;
		if (s0_clk_en)
			s1_req_signed <= io_cpu_req_bits_signed;
		if (s0_clk_en)
			s1_req_dprv <= io_cpu_req_bits_dprv;
		if (s0_clk_en)
			s1_tlb_req_vaddr <= s0_req_addr;
		if (s0_clk_en)
			s1_tlb_req_size <= io_cpu_req_bits_size;
		if (s0_clk_en)
			s1_tlb_req_cmd <= io_cpu_req_bits_cmd;
		if (s0_clk_en)
			s1_tlb_req_prv <= io_cpu_req_bits_dprv;
		s1_flush_valid <= (_s1_flush_valid_T & ~s1_flush_valid) & _s2_cannot_victimize_T;
		if (reset)
			uncachedInFlight_0 <= 1'h0;
		else if (_T_261) begin
			if (grantIsCached)
				uncachedInFlight_0 <= _GEN_158;
			else if (d_last)
				uncachedInFlight_0 <= 1'h0;
			else
				uncachedInFlight_0 <= _GEN_158;
		end
		else
			uncachedInFlight_0 <= _GEN_158;
		if (_T_244)
			uncachedReqs_0_addr <= s2_req_addr;
		if (_T_244)
			uncachedReqs_0_tag <= s2_req_tag;
		if (_T_244)
			uncachedReqs_0_size <= s2_req_size;
		if (_T_244)
			uncachedReqs_0_signed <= s2_req_signed;
		if (s0_clk_en)
			s1_did_read <= _s1_did_read_T_54;
		if (s0_clk_en)
			s1_read_mask <= dataArb_io_in_3_bits_wordMask;
		if (_T_261) begin
			if (grantIsCached)
				s2_req_addr <= _GEN_40;
			else if (data_1)
				s2_req_addr <= _s2_req_addr_T_1;
			else
				s2_req_addr <= _GEN_40;
		end
		else
			s2_req_addr <= _GEN_40;
		if (_T_261) begin
			if (grantIsCached)
				s2_req_tag <= _GEN_41;
			else if (data_1)
				s2_req_tag <= uncachedReqs_0_tag;
			else
				s2_req_tag <= _GEN_41;
		end
		else
			s2_req_tag <= _GEN_41;
		if (_T_261) begin
			if (grantIsCached)
				s2_req_size <= _GEN_43;
			else if (data_1)
				s2_req_size <= uncachedReqs_0_size;
			else
				s2_req_size <= _GEN_43;
		end
		else
			s2_req_size <= _GEN_43;
		if (_T_261) begin
			if (grantIsCached)
				s2_req_signed <= _GEN_44;
			else if (data_1)
				s2_req_signed <= uncachedReqs_0_signed;
			else
				s2_req_signed <= _GEN_44;
		end
		else
			s2_req_signed <= _GEN_44;
		if (s1_valid_not_nacked | s1_flush_valid)
			s2_req_dprv <= s1_req_dprv;
		if (s1_valid_not_nacked | s1_flush_valid)
			s2_req_no_xcpt <= s1_req_no_xcpt;
		if (s1_valid_not_nacked | s1_flush_valid)
			s2_tlb_xcpt_pf_ld <= tlb_io_resp_pf_ld;
		if (s1_valid_not_nacked | s1_flush_valid)
			s2_tlb_xcpt_pf_st <= tlb_io_resp_pf_st;
		if (s1_valid_not_nacked | s1_flush_valid)
			s2_tlb_xcpt_ae_ld <= tlb_io_resp_ae_ld;
		if (s1_valid_not_nacked | s1_flush_valid)
			s2_tlb_xcpt_ae_st <= tlb_io_resp_ae_st;
		if (s1_valid_not_nacked | s1_flush_valid)
			s2_tlb_xcpt_ma_ld <= tlb_io_resp_ma_ld;
		if (s1_valid_not_nacked | s1_flush_valid)
			s2_tlb_xcpt_ma_st <= tlb_io_resp_ma_st;
		if (_T_261)
			if (!grantIsCached)
				if (data_1)
					s2_uncached_resp_addr <= uncachedReqs_0_addr;
		if (_T_34)
			s2_vaddr_r <= s1_vaddr;
		s2_flush_valid_pre_tag_ecc <= s1_flush_valid;
		if (data_1 & (blockUncachedGrant | s1_valid)) begin
			if (auto_out_d_valid)
				blockUncachedGrant <= _T_284;
			else
				blockUncachedGrant <= dataArb_io_out_valid;
		end
		else
			blockUncachedGrant <= dataArb_io_out_valid;
		if (reset)
			counter <= 10'h000;
		else if (_T_261)
			if (d_first) begin
				if (beats1_opdata)
					counter <= beats1_decode;
				else
					counter <= 10'h000;
			end
			else
				counter <= counter1;
		if (en)
			s2_data <= _s2_data_T_6;
		if (_pstore1_cmd_T)
			pstore1_cmd <= s1_req_cmd;
		if (_pstore1_cmd_T)
			pstore1_data <= io_cpu_s1_data_data;
		if (_pstore1_cmd_T)
			pstore1_rmw_r <= _pstore1_rmw_T_52;
		pstore_drain_on_miss_REG <= io_cpu_s2_nack;
		if (advance_pstore1)
			pstore2_storegen_data_r <= pstore1_storegen_data[7:0];
		if (advance_pstore1)
			pstore2_storegen_data_r_1 <= pstore1_storegen_data[15:8];
		if (advance_pstore1)
			pstore2_storegen_data_r_2 <= pstore1_storegen_data[23:16];
		if (advance_pstore1)
			pstore2_storegen_data_r_3 <= pstore1_storegen_data[31:24];
		io_cpu_s2_xcpt_REG <= (tlb_io_req_valid & _io_cpu_ordered_T) & _s1_valid_not_nacked_T;
		doUncachedResp <= io_cpu_replay_next;
	end
endmodule
module ICache (
	clock,
	reset,
	auto_master_out_a_ready,
	auto_master_out_a_valid,
	auto_master_out_a_bits_address,
	auto_master_out_d_valid,
	auto_master_out_d_bits_opcode,
	auto_master_out_d_bits_size,
	auto_master_out_d_bits_data,
	auto_master_out_d_bits_corrupt,
	io_req_ready,
	io_req_valid,
	io_req_bits_addr,
	io_s1_paddr,
	io_s1_kill,
	io_s2_kill,
	io_resp_valid,
	io_resp_bits_data,
	io_resp_bits_ae,
	io_invalidate
);
	input clock;
	input reset;
	input auto_master_out_a_ready;
	output wire auto_master_out_a_valid;
	output wire [31:0] auto_master_out_a_bits_address;
	input auto_master_out_d_valid;
	input [2:0] auto_master_out_d_bits_opcode;
	input [3:0] auto_master_out_d_bits_size;
	input [31:0] auto_master_out_d_bits_data;
	input auto_master_out_d_bits_corrupt;
	output wire io_req_ready;
	input io_req_valid;
	input [31:0] io_req_bits_addr;
	input [31:0] io_s1_paddr;
	input io_s1_kill;
	input io_s2_kill;
	output wire io_resp_valid;
	output wire [31:0] io_resp_bits_data;
	output wire io_resp_bits_ae;
	input io_invalidate;
	wire [5:0] tag_array_RW0_addr;
	wire tag_array_RW0_en;
	wire tag_array_RW0_clk;
	wire tag_array_RW0_wmode;
	wire [20:0] tag_array_RW0_wdata_0;
	wire [20:0] tag_array_RW0_rdata_0;
	wire [9:0] data_arrays_0_RW0_addr;
	wire data_arrays_0_RW0_en;
	wire data_arrays_0_RW0_clk;
	wire data_arrays_0_RW0_wmode;
	wire [31:0] data_arrays_0_RW0_wdata_0;
	wire [31:0] data_arrays_0_RW0_rdata_0;
	wire s0_valid = io_req_ready & io_req_valid;
	reg s1_valid;
	reg [63:0] vb_array;
	wire [5:0] s1_idx = io_s1_paddr[11:6];
	wire [6:0] _s1_vb_T = {1'h0, s1_idx};
	wire [63:0] _s1_vb_T_1 = vb_array >> _s1_vb_T;
	wire s1_vb = _s1_vb_T_1[0];
	wire [19:0] tag = tag_array_RW0_rdata_0[19:0];
	wire [19:0] s1_tag = io_s1_paddr[31:12];
	wire tagMatch = s1_vb & (tag == s1_tag);
	wire _s1_tag_hit_0_T = tagMatch;
	wire s1_hit = tagMatch;
	reg s2_valid;
	reg s2_hit;
	reg invalidated;
	reg refill_valid;
	wire s2_miss = (s2_valid & ~s2_hit) & ~io_s2_kill;
	reg s2_request_refill_REG;
	wire s2_request_refill = s2_miss & s2_request_refill_REG;
	wire refill_fire = auto_master_out_a_ready & s2_request_refill;
	wire s1_can_request_refill = ~(s2_miss | refill_valid);
	wire _refill_paddr_T = s1_valid & s1_can_request_refill;
	reg [31:0] refill_paddr;
	wire [19:0] refill_tag = refill_paddr[31:12];
	wire [5:0] refill_idx = refill_paddr[11:6];
	wire refill_one_beat_opdata = auto_master_out_d_bits_opcode[0];
	wire refill_one_beat = auto_master_out_d_valid & refill_one_beat_opdata;
	wire [26:0] _beats1_decode_T_1 = 27'h0000fff << auto_master_out_d_bits_size;
	wire [11:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[11:0];
	wire [9:0] beats1_decode = _beats1_decode_T_3[11:2];
	wire [9:0] beats1 = (refill_one_beat_opdata ? beats1_decode : 10'h000);
	reg [9:0] counter;
	wire [9:0] counter1 = counter - 10'h001;
	wire first = counter == 10'h000;
	wire last = (counter == 10'h001) | (beats1 == 10'h000);
	wire d_done = last & auto_master_out_d_valid;
	wire [9:0] _count_T = ~counter1;
	wire [9:0] refill_cnt = beats1 & _count_T;
	wire refill_done = refill_one_beat & d_done;
	wire _tag_rdata_T_2 = ~refill_done & s0_valid;
	reg accruedRefillError;
	wire refillError = auto_master_out_d_bits_corrupt | ((refill_cnt > 10'h000) & accruedRefillError);
	wire [6:0] _vb_array_T = {1'h0, refill_idx};
	wire _vb_array_T_1 = ~invalidated;
	wire [127:0] _vb_array_T_3 = 128'h00000000000000000000000000000001 << _vb_array_T;
	wire [127:0] _GEN_40 = {64'd0, vb_array};
	wire [127:0] _vb_array_T_4 = _GEN_40 | _vb_array_T_3;
	wire [63:0] _vb_array_T_5 = ~vb_array;
	wire [127:0] _GEN_41 = {64'd0, _vb_array_T_5};
	wire [127:0] _vb_array_T_6 = _GEN_41 | _vb_array_T_3;
	wire [127:0] _vb_array_T_7 = ~_vb_array_T_6;
	wire [127:0] _vb_array_T_8 = (refill_done & ~invalidated ? _vb_array_T_4 : _vb_array_T_7);
	wire [127:0] _GEN_16 = (refill_one_beat ? _vb_array_T_8 : {64'd0, vb_array});
	wire [127:0] _GEN_17 = (io_invalidate ? 128'h00000000000000000000000000000000 : _GEN_16);
	wire _GEN_18 = io_invalidate | invalidated;
	wire tl_error = tag_array_RW0_rdata_0[20];
	wire s1_tl_error_0 = tagMatch & tl_error;
	wire wen = refill_one_beat & _vb_array_T_1;
	wire [9:0] _mem_idx_T = {refill_idx, 4'h0};
	wire [9:0] _mem_idx_T_1 = _mem_idx_T | refill_cnt;
	wire _dout_T_1 = ~wen & s0_valid;
	wire [31:0] s1_dout_0 = data_arrays_0_RW0_rdata_0;
	reg [31:0] s2_dout_0;
	wire _s2_tl_error_T = |s1_tl_error_0;
	reg s2_tl_error;
	wire _GEN_38 = refill_fire | refill_valid;
	tag_array tag_array(
		.RW0_addr(tag_array_RW0_addr),
		.RW0_en(tag_array_RW0_en),
		.RW0_clk(tag_array_RW0_clk),
		.RW0_wmode(tag_array_RW0_wmode),
		.RW0_wdata_0(tag_array_RW0_wdata_0),
		.RW0_rdata_0(tag_array_RW0_rdata_0)
	);
	data_arrays_0_0 data_arrays_0(
		.RW0_addr(data_arrays_0_RW0_addr),
		.RW0_en(data_arrays_0_RW0_en),
		.RW0_clk(data_arrays_0_RW0_clk),
		.RW0_wmode(data_arrays_0_RW0_wmode),
		.RW0_wdata_0(data_arrays_0_RW0_wdata_0),
		.RW0_rdata_0(data_arrays_0_RW0_rdata_0)
	);
	assign auto_master_out_a_valid = s2_miss & s2_request_refill_REG;
	assign auto_master_out_a_bits_address = {refill_paddr[31:6], 6'h00};
	assign io_req_ready = ~refill_one_beat;
	assign io_resp_valid = s2_valid & s2_hit;
	assign io_resp_bits_data = s2_dout_0;
	assign io_resp_bits_ae = s2_tl_error;
	assign tag_array_RW0_clk = clock;
	assign tag_array_RW0_wdata_0 = {refillError, refill_tag};
	assign data_arrays_0_RW0_clk = clock;
	assign data_arrays_0_RW0_wdata_0 = auto_master_out_d_bits_data;
	assign tag_array_RW0_en = _tag_rdata_T_2 | refill_done;
	assign tag_array_RW0_wmode = refill_one_beat & d_done;
	assign tag_array_RW0_addr = (refill_done ? refill_idx : io_req_bits_addr[11:6]);
	assign data_arrays_0_RW0_en = _dout_T_1 | wen;
	assign data_arrays_0_RW0_wmode = refill_one_beat & _vb_array_T_1;
	assign data_arrays_0_RW0_addr = (refill_one_beat ? _mem_idx_T_1 : io_req_bits_addr[11:2]);
	always @(posedge clock) begin
		if (reset)
			s1_valid <= 1'h0;
		else
			s1_valid <= s0_valid;
		if (reset)
			vb_array <= 64'h0000000000000000;
		else
			vb_array <= _GEN_17[63:0];
		if (reset)
			s2_valid <= 1'h0;
		else
			s2_valid <= s1_valid & ~io_s1_kill;
		s2_hit <= _s1_tag_hit_0_T;
		if (~refill_valid)
			invalidated <= 1'h0;
		else
			invalidated <= _GEN_18;
		if (reset)
			refill_valid <= 1'h0;
		else if (refill_done)
			refill_valid <= 1'h0;
		else
			refill_valid <= _GEN_38;
		s2_request_refill_REG <= ~(s2_miss | refill_valid);
		if (_refill_paddr_T)
			refill_paddr <= io_s1_paddr;
		if (reset)
			counter <= 10'h000;
		else if (auto_master_out_d_valid)
			if (first) begin
				if (refill_one_beat_opdata)
					counter <= beats1_decode;
				else
					counter <= 10'h000;
			end
			else
				counter <= counter1;
		if (refill_one_beat)
			accruedRefillError <= refillError;
		if (s1_valid)
			s2_dout_0 <= s1_dout_0;
		if (s1_valid)
			s2_tl_error <= _s2_tl_error_T;
	end
endmodule
module ShiftQueue (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_pc,
	io_enq_bits_data,
	io_enq_bits_xcpt_ae_inst,
	io_enq_bits_replay,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_pc,
	io_deq_bits_data,
	io_deq_bits_xcpt_ae_inst,
	io_deq_bits_replay,
	io_mask
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [31:0] io_enq_bits_pc;
	input [31:0] io_enq_bits_data;
	input io_enq_bits_xcpt_ae_inst;
	input io_enq_bits_replay;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [31:0] io_deq_bits_pc;
	output wire [31:0] io_deq_bits_data;
	output wire io_deq_bits_xcpt_ae_inst;
	output wire io_deq_bits_replay;
	output wire [4:0] io_mask;
	reg valid_0;
	reg valid_1;
	reg valid_2;
	reg valid_3;
	reg valid_4;
	reg [31:0] elts_0_pc;
	reg [31:0] elts_0_data;
	reg elts_0_xcpt_ae_inst;
	reg elts_0_replay;
	reg [31:0] elts_1_pc;
	reg [31:0] elts_1_data;
	reg elts_1_xcpt_ae_inst;
	reg elts_1_replay;
	reg [31:0] elts_2_pc;
	reg [31:0] elts_2_data;
	reg elts_2_xcpt_ae_inst;
	reg elts_2_replay;
	reg [31:0] elts_3_pc;
	reg [31:0] elts_3_data;
	reg elts_3_xcpt_ae_inst;
	reg elts_3_replay;
	reg [31:0] elts_4_pc;
	reg [31:0] elts_4_data;
	reg elts_4_xcpt_ae_inst;
	reg elts_4_replay;
	wire _wen_T = io_enq_ready & io_enq_valid;
	wire _wen_T_2 = _wen_T & valid_0;
	wire _wen_T_3 = valid_1 | (_wen_T & valid_0);
	wire _wen_T_6 = ~valid_0;
	wire _wen_T_7 = _wen_T & ~valid_0;
	wire wen = (io_deq_ready ? _wen_T_3 : _wen_T_7);
	wire _valid_0_T_6 = _wen_T | valid_0;
	wire _wen_T_10 = _wen_T & valid_1;
	wire _wen_T_11 = valid_2 | (_wen_T & valid_1);
	wire _wen_T_15 = _wen_T_2 & ~valid_1;
	wire wen_1 = (io_deq_ready ? _wen_T_11 : _wen_T_15);
	wire _valid_1_T_6 = _wen_T_2 | valid_1;
	wire _wen_T_18 = _wen_T & valid_2;
	wire _wen_T_19 = valid_3 | (_wen_T & valid_2);
	wire _wen_T_23 = _wen_T_10 & ~valid_2;
	wire wen_2 = (io_deq_ready ? _wen_T_19 : _wen_T_23);
	wire _valid_2_T_6 = _wen_T_10 | valid_2;
	wire _wen_T_26 = _wen_T & valid_3;
	wire _wen_T_27 = valid_4 | (_wen_T & valid_3);
	wire _wen_T_31 = _wen_T_18 & ~valid_3;
	wire wen_3 = (io_deq_ready ? _wen_T_27 : _wen_T_31);
	wire _valid_3_T_6 = _wen_T_18 | valid_3;
	wire _wen_T_34 = _wen_T & valid_4;
	wire _wen_T_39 = _wen_T_26 & ~valid_4;
	wire wen_4 = (io_deq_ready ? _wen_T_34 : _wen_T_39);
	wire _valid_4_T_6 = _wen_T_26 | valid_4;
	wire [1:0] io_mask_lo = {valid_1, valid_0};
	wire [2:0] io_mask_hi = {valid_4, valid_3, valid_2};
	assign io_enq_ready = ~valid_4;
	assign io_deq_valid = io_enq_valid | valid_0;
	assign io_deq_bits_pc = (_wen_T_6 ? io_enq_bits_pc : elts_0_pc);
	assign io_deq_bits_data = (_wen_T_6 ? io_enq_bits_data : elts_0_data);
	assign io_deq_bits_xcpt_ae_inst = (_wen_T_6 ? io_enq_bits_xcpt_ae_inst : elts_0_xcpt_ae_inst);
	assign io_deq_bits_replay = (_wen_T_6 ? io_enq_bits_replay : elts_0_replay);
	assign io_mask = {io_mask_hi, io_mask_lo};
	always @(posedge clock) begin
		if (reset)
			valid_0 <= 1'h0;
		else if (io_deq_ready)
			valid_0 <= _wen_T_3;
		else
			valid_0 <= _valid_0_T_6;
		if (reset)
			valid_1 <= 1'h0;
		else if (io_deq_ready)
			valid_1 <= _wen_T_11;
		else
			valid_1 <= _valid_1_T_6;
		if (reset)
			valid_2 <= 1'h0;
		else if (io_deq_ready)
			valid_2 <= _wen_T_19;
		else
			valid_2 <= _valid_2_T_6;
		if (reset)
			valid_3 <= 1'h0;
		else if (io_deq_ready)
			valid_3 <= _wen_T_27;
		else
			valid_3 <= _valid_3_T_6;
		if (reset)
			valid_4 <= 1'h0;
		else if (io_deq_ready)
			valid_4 <= _wen_T_34;
		else
			valid_4 <= _valid_4_T_6;
		if (wen)
			if (valid_1)
				elts_0_pc <= elts_1_pc;
			else
				elts_0_pc <= io_enq_bits_pc;
		if (wen)
			if (valid_1)
				elts_0_data <= elts_1_data;
			else
				elts_0_data <= io_enq_bits_data;
		if (wen)
			if (valid_1)
				elts_0_xcpt_ae_inst <= elts_1_xcpt_ae_inst;
			else
				elts_0_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
		if (wen)
			if (valid_1)
				elts_0_replay <= elts_1_replay;
			else
				elts_0_replay <= io_enq_bits_replay;
		if (wen_1)
			if (valid_2)
				elts_1_pc <= elts_2_pc;
			else
				elts_1_pc <= io_enq_bits_pc;
		if (wen_1)
			if (valid_2)
				elts_1_data <= elts_2_data;
			else
				elts_1_data <= io_enq_bits_data;
		if (wen_1)
			if (valid_2)
				elts_1_xcpt_ae_inst <= elts_2_xcpt_ae_inst;
			else
				elts_1_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
		if (wen_1)
			if (valid_2)
				elts_1_replay <= elts_2_replay;
			else
				elts_1_replay <= io_enq_bits_replay;
		if (wen_2)
			if (valid_3)
				elts_2_pc <= elts_3_pc;
			else
				elts_2_pc <= io_enq_bits_pc;
		if (wen_2)
			if (valid_3)
				elts_2_data <= elts_3_data;
			else
				elts_2_data <= io_enq_bits_data;
		if (wen_2)
			if (valid_3)
				elts_2_xcpt_ae_inst <= elts_3_xcpt_ae_inst;
			else
				elts_2_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
		if (wen_2)
			if (valid_3)
				elts_2_replay <= elts_3_replay;
			else
				elts_2_replay <= io_enq_bits_replay;
		if (wen_3)
			if (valid_4)
				elts_3_pc <= elts_4_pc;
			else
				elts_3_pc <= io_enq_bits_pc;
		if (wen_3)
			if (valid_4)
				elts_3_data <= elts_4_data;
			else
				elts_3_data <= io_enq_bits_data;
		if (wen_3)
			if (valid_4)
				elts_3_xcpt_ae_inst <= elts_4_xcpt_ae_inst;
			else
				elts_3_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
		if (wen_3)
			if (valid_4)
				elts_3_replay <= elts_4_replay;
			else
				elts_3_replay <= io_enq_bits_replay;
		if (wen_4)
			elts_4_pc <= io_enq_bits_pc;
		if (wen_4)
			elts_4_data <= io_enq_bits_data;
		if (wen_4)
			elts_4_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
		if (wen_4)
			elts_4_replay <= io_enq_bits_replay;
	end
endmodule
module TLB_1 (
	io_req_bits_vaddr,
	io_resp_paddr,
	io_resp_ae_inst,
	io_ptw_status_debug,
	io_ptw_pmp_0_cfg_l,
	io_ptw_pmp_0_cfg_a,
	io_ptw_pmp_0_cfg_x,
	io_ptw_pmp_0_cfg_w,
	io_ptw_pmp_0_cfg_r,
	io_ptw_pmp_0_addr,
	io_ptw_pmp_0_mask,
	io_ptw_pmp_1_cfg_l,
	io_ptw_pmp_1_cfg_a,
	io_ptw_pmp_1_cfg_x,
	io_ptw_pmp_1_cfg_w,
	io_ptw_pmp_1_cfg_r,
	io_ptw_pmp_1_addr,
	io_ptw_pmp_1_mask,
	io_ptw_pmp_2_cfg_l,
	io_ptw_pmp_2_cfg_a,
	io_ptw_pmp_2_cfg_x,
	io_ptw_pmp_2_cfg_w,
	io_ptw_pmp_2_cfg_r,
	io_ptw_pmp_2_addr,
	io_ptw_pmp_2_mask,
	io_ptw_pmp_3_cfg_l,
	io_ptw_pmp_3_cfg_a,
	io_ptw_pmp_3_cfg_x,
	io_ptw_pmp_3_cfg_w,
	io_ptw_pmp_3_cfg_r,
	io_ptw_pmp_3_addr,
	io_ptw_pmp_3_mask,
	io_ptw_pmp_4_cfg_l,
	io_ptw_pmp_4_cfg_a,
	io_ptw_pmp_4_cfg_x,
	io_ptw_pmp_4_cfg_w,
	io_ptw_pmp_4_cfg_r,
	io_ptw_pmp_4_addr,
	io_ptw_pmp_4_mask,
	io_ptw_pmp_5_cfg_l,
	io_ptw_pmp_5_cfg_a,
	io_ptw_pmp_5_cfg_x,
	io_ptw_pmp_5_cfg_w,
	io_ptw_pmp_5_cfg_r,
	io_ptw_pmp_5_addr,
	io_ptw_pmp_5_mask,
	io_ptw_pmp_6_cfg_l,
	io_ptw_pmp_6_cfg_a,
	io_ptw_pmp_6_cfg_x,
	io_ptw_pmp_6_cfg_w,
	io_ptw_pmp_6_cfg_r,
	io_ptw_pmp_6_addr,
	io_ptw_pmp_6_mask,
	io_ptw_pmp_7_cfg_l,
	io_ptw_pmp_7_cfg_a,
	io_ptw_pmp_7_cfg_x,
	io_ptw_pmp_7_cfg_w,
	io_ptw_pmp_7_cfg_r,
	io_ptw_pmp_7_addr,
	io_ptw_pmp_7_mask
);
	input [31:0] io_req_bits_vaddr;
	output wire [31:0] io_resp_paddr;
	output wire io_resp_ae_inst;
	input io_ptw_status_debug;
	input io_ptw_pmp_0_cfg_l;
	input [1:0] io_ptw_pmp_0_cfg_a;
	input io_ptw_pmp_0_cfg_x;
	input io_ptw_pmp_0_cfg_w;
	input io_ptw_pmp_0_cfg_r;
	input [29:0] io_ptw_pmp_0_addr;
	input [31:0] io_ptw_pmp_0_mask;
	input io_ptw_pmp_1_cfg_l;
	input [1:0] io_ptw_pmp_1_cfg_a;
	input io_ptw_pmp_1_cfg_x;
	input io_ptw_pmp_1_cfg_w;
	input io_ptw_pmp_1_cfg_r;
	input [29:0] io_ptw_pmp_1_addr;
	input [31:0] io_ptw_pmp_1_mask;
	input io_ptw_pmp_2_cfg_l;
	input [1:0] io_ptw_pmp_2_cfg_a;
	input io_ptw_pmp_2_cfg_x;
	input io_ptw_pmp_2_cfg_w;
	input io_ptw_pmp_2_cfg_r;
	input [29:0] io_ptw_pmp_2_addr;
	input [31:0] io_ptw_pmp_2_mask;
	input io_ptw_pmp_3_cfg_l;
	input [1:0] io_ptw_pmp_3_cfg_a;
	input io_ptw_pmp_3_cfg_x;
	input io_ptw_pmp_3_cfg_w;
	input io_ptw_pmp_3_cfg_r;
	input [29:0] io_ptw_pmp_3_addr;
	input [31:0] io_ptw_pmp_3_mask;
	input io_ptw_pmp_4_cfg_l;
	input [1:0] io_ptw_pmp_4_cfg_a;
	input io_ptw_pmp_4_cfg_x;
	input io_ptw_pmp_4_cfg_w;
	input io_ptw_pmp_4_cfg_r;
	input [29:0] io_ptw_pmp_4_addr;
	input [31:0] io_ptw_pmp_4_mask;
	input io_ptw_pmp_5_cfg_l;
	input [1:0] io_ptw_pmp_5_cfg_a;
	input io_ptw_pmp_5_cfg_x;
	input io_ptw_pmp_5_cfg_w;
	input io_ptw_pmp_5_cfg_r;
	input [29:0] io_ptw_pmp_5_addr;
	input [31:0] io_ptw_pmp_5_mask;
	input io_ptw_pmp_6_cfg_l;
	input [1:0] io_ptw_pmp_6_cfg_a;
	input io_ptw_pmp_6_cfg_x;
	input io_ptw_pmp_6_cfg_w;
	input io_ptw_pmp_6_cfg_r;
	input [29:0] io_ptw_pmp_6_addr;
	input [31:0] io_ptw_pmp_6_mask;
	input io_ptw_pmp_7_cfg_l;
	input [1:0] io_ptw_pmp_7_cfg_a;
	input io_ptw_pmp_7_cfg_x;
	input io_ptw_pmp_7_cfg_w;
	input io_ptw_pmp_7_cfg_r;
	input [29:0] io_ptw_pmp_7_addr;
	input [31:0] io_ptw_pmp_7_mask;
	wire [1:0] pmp_io_prv;
	wire pmp_io_pmp_0_cfg_l;
	wire [1:0] pmp_io_pmp_0_cfg_a;
	wire pmp_io_pmp_0_cfg_x;
	wire pmp_io_pmp_0_cfg_w;
	wire pmp_io_pmp_0_cfg_r;
	wire [29:0] pmp_io_pmp_0_addr;
	wire [31:0] pmp_io_pmp_0_mask;
	wire pmp_io_pmp_1_cfg_l;
	wire [1:0] pmp_io_pmp_1_cfg_a;
	wire pmp_io_pmp_1_cfg_x;
	wire pmp_io_pmp_1_cfg_w;
	wire pmp_io_pmp_1_cfg_r;
	wire [29:0] pmp_io_pmp_1_addr;
	wire [31:0] pmp_io_pmp_1_mask;
	wire pmp_io_pmp_2_cfg_l;
	wire [1:0] pmp_io_pmp_2_cfg_a;
	wire pmp_io_pmp_2_cfg_x;
	wire pmp_io_pmp_2_cfg_w;
	wire pmp_io_pmp_2_cfg_r;
	wire [29:0] pmp_io_pmp_2_addr;
	wire [31:0] pmp_io_pmp_2_mask;
	wire pmp_io_pmp_3_cfg_l;
	wire [1:0] pmp_io_pmp_3_cfg_a;
	wire pmp_io_pmp_3_cfg_x;
	wire pmp_io_pmp_3_cfg_w;
	wire pmp_io_pmp_3_cfg_r;
	wire [29:0] pmp_io_pmp_3_addr;
	wire [31:0] pmp_io_pmp_3_mask;
	wire pmp_io_pmp_4_cfg_l;
	wire [1:0] pmp_io_pmp_4_cfg_a;
	wire pmp_io_pmp_4_cfg_x;
	wire pmp_io_pmp_4_cfg_w;
	wire pmp_io_pmp_4_cfg_r;
	wire [29:0] pmp_io_pmp_4_addr;
	wire [31:0] pmp_io_pmp_4_mask;
	wire pmp_io_pmp_5_cfg_l;
	wire [1:0] pmp_io_pmp_5_cfg_a;
	wire pmp_io_pmp_5_cfg_x;
	wire pmp_io_pmp_5_cfg_w;
	wire pmp_io_pmp_5_cfg_r;
	wire [29:0] pmp_io_pmp_5_addr;
	wire [31:0] pmp_io_pmp_5_mask;
	wire pmp_io_pmp_6_cfg_l;
	wire [1:0] pmp_io_pmp_6_cfg_a;
	wire pmp_io_pmp_6_cfg_x;
	wire pmp_io_pmp_6_cfg_w;
	wire pmp_io_pmp_6_cfg_r;
	wire [29:0] pmp_io_pmp_6_addr;
	wire [31:0] pmp_io_pmp_6_mask;
	wire pmp_io_pmp_7_cfg_l;
	wire [1:0] pmp_io_pmp_7_cfg_a;
	wire pmp_io_pmp_7_cfg_x;
	wire pmp_io_pmp_7_cfg_w;
	wire pmp_io_pmp_7_cfg_r;
	wire [29:0] pmp_io_pmp_7_addr;
	wire [31:0] pmp_io_pmp_7_mask;
	wire [31:0] pmp_io_addr;
	wire pmp_io_r;
	wire pmp_io_w;
	wire pmp_io_x;
	wire [19:0] vpn = io_req_bits_vaddr[31:12];
	wire [19:0] mpu_ppn = io_req_bits_vaddr[31:12];
	wire [31:0] mpu_physaddr = {mpu_ppn, io_req_bits_vaddr[11:0]};
	wire [2:0] mpu_priv = {io_ptw_status_debug, 2'h3};
	wire [31:0] _legal_address_T = mpu_physaddr ^ 32'h00003000;
	wire [32:0] _legal_address_T_1 = {1'b0, $signed(_legal_address_T)};
	wire [32:0] _legal_address_T_3 = $signed(_legal_address_T_1) & -33'sh000001000;
	wire _legal_address_T_4 = $signed(_legal_address_T_3) == 33'sh000000000;
	wire [31:0] _legal_address_T_5 = mpu_physaddr ^ 32'h00004000;
	wire [32:0] _legal_address_T_6 = {1'b0, $signed(_legal_address_T_5)};
	wire [32:0] _legal_address_T_8 = $signed(_legal_address_T_6) & -33'sh000001000;
	wire _legal_address_T_9 = $signed(_legal_address_T_8) == 33'sh000000000;
	wire [31:0] _legal_address_T_10 = mpu_physaddr ^ 32'h10000000;
	wire [32:0] _legal_address_T_11 = {1'b0, $signed(_legal_address_T_10)};
	wire [32:0] _legal_address_T_13 = $signed(_legal_address_T_11) & -33'sh000001000;
	wire _legal_address_T_14 = $signed(_legal_address_T_13) == 33'sh000000000;
	wire [31:0] _legal_address_T_15 = mpu_physaddr ^ 32'h00020000;
	wire [32:0] _legal_address_T_16 = {1'b0, $signed(_legal_address_T_15)};
	wire [32:0] _legal_address_T_18 = $signed(_legal_address_T_16) & -33'sh000010000;
	wire _legal_address_T_19 = $signed(_legal_address_T_18) == 33'sh000000000;
	wire [31:0] _legal_address_T_20 = mpu_physaddr ^ 32'h54000000;
	wire [32:0] _legal_address_T_21 = {1'b0, $signed(_legal_address_T_20)};
	wire [32:0] _legal_address_T_23 = $signed(_legal_address_T_21) & -33'sh000001000;
	wire _legal_address_T_24 = $signed(_legal_address_T_23) == 33'sh000000000;
	wire [31:0] _legal_address_T_25 = mpu_physaddr ^ 32'h0c000000;
	wire [32:0] _legal_address_T_26 = {1'b0, $signed(_legal_address_T_25)};
	wire [32:0] _legal_address_T_28 = $signed(_legal_address_T_26) & -33'sh004000000;
	wire _legal_address_T_29 = $signed(_legal_address_T_28) == 33'sh000000000;
	wire [31:0] _legal_address_T_30 = mpu_physaddr ^ 32'h02000000;
	wire [32:0] _legal_address_T_31 = {1'b0, $signed(_legal_address_T_30)};
	wire [32:0] _legal_address_T_33 = $signed(_legal_address_T_31) & -33'sh000010000;
	wire _legal_address_T_34 = $signed(_legal_address_T_33) == 33'sh000000000;
	wire [32:0] _legal_address_T_36 = {1'b0, $signed(mpu_physaddr)};
	wire [32:0] _legal_address_T_38 = $signed(_legal_address_T_36) & -33'sh000001000;
	wire _legal_address_T_39 = $signed(_legal_address_T_38) == 33'sh000000000;
	wire [31:0] _legal_address_T_40 = mpu_physaddr ^ 32'h80000000;
	wire [32:0] _legal_address_T_41 = {1'b0, $signed(_legal_address_T_40)};
	wire [32:0] _legal_address_T_43 = $signed(_legal_address_T_41) & -33'sh000004000;
	wire _legal_address_T_44 = $signed(_legal_address_T_43) == 33'sh000000000;
	wire [31:0] _legal_address_T_45 = mpu_physaddr ^ 32'h00010000;
	wire [32:0] _legal_address_T_46 = {1'b0, $signed(_legal_address_T_45)};
	wire [32:0] _legal_address_T_48 = $signed(_legal_address_T_46) & -33'sh000010000;
	wire _legal_address_T_49 = $signed(_legal_address_T_48) == 33'sh000000000;
	wire [31:0] _legal_address_T_50 = mpu_physaddr ^ 32'h00100000;
	wire [32:0] _legal_address_T_51 = {1'b0, $signed(_legal_address_T_50)};
	wire [32:0] _legal_address_T_53 = $signed(_legal_address_T_51) & -33'sh000001000;
	wire _legal_address_T_54 = $signed(_legal_address_T_53) == 33'sh000000000;
	wire [31:0] _legal_address_T_55 = mpu_physaddr ^ 32'h00110000;
	wire [32:0] _legal_address_T_56 = {1'b0, $signed(_legal_address_T_55)};
	wire [32:0] _legal_address_T_58 = $signed(_legal_address_T_56) & -33'sh000001000;
	wire _legal_address_T_59 = $signed(_legal_address_T_58) == 33'sh000000000;
	wire legal_address = ((((((((((_legal_address_T_4 | _legal_address_T_9) | _legal_address_T_14) | _legal_address_T_19) | _legal_address_T_24) | _legal_address_T_29) | _legal_address_T_34) | _legal_address_T_39) | _legal_address_T_44) | _legal_address_T_49) | _legal_address_T_54) | _legal_address_T_59;
	wire [32:0] _homogeneous_T_76 = $signed(_legal_address_T_36) & 33'sh016134000;
	wire _homogeneous_T_77 = $signed(_homogeneous_T_76) == 33'sh000000000;
	wire [32:0] _homogeneous_T_81 = $signed(_legal_address_T_46) & 33'sh096130000;
	wire _homogeneous_T_82 = $signed(_homogeneous_T_81) == 33'sh000000000;
	wire [32:0] _homogeneous_T_86 = $signed(_legal_address_T_16) & 33'sh096130000;
	wire _homogeneous_T_87 = $signed(_homogeneous_T_86) == 33'sh000000000;
	wire [32:0] _homogeneous_T_91 = $signed(_legal_address_T_11) & 33'sh096136000;
	wire _homogeneous_T_92 = $signed(_homogeneous_T_91) == 33'sh000000000;
	wire _homogeneous_T_96 = ((_homogeneous_T_77 | _homogeneous_T_82) | _homogeneous_T_87) | _homogeneous_T_92;
	wire deny_access_to_debug = (mpu_priv <= 3'h3) & _legal_address_T_39;
	wire _prot_r_T_6 = ~deny_access_to_debug;
	wire _prot_x_T_55 = legal_address & _homogeneous_T_96;
	wire prot_x = (_prot_x_T_55 & _prot_r_T_6) & pmp_io_x;
	wire [1:0] _px_array_T_1 = (prot_x ? 2'h3 : 2'h0);
	wire [6:0] px_array = {_px_array_T_1, 5'h00};
	wire [6:0] _io_resp_ae_inst_T = ~px_array;
	wire [6:0] _io_resp_ae_inst_T_1 = _io_resp_ae_inst_T & 7'h40;
	PMPChecker pmp(
		.io_prv(pmp_io_prv),
		.io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
		.io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
		.io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
		.io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
		.io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
		.io_pmp_0_addr(pmp_io_pmp_0_addr),
		.io_pmp_0_mask(pmp_io_pmp_0_mask),
		.io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
		.io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
		.io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
		.io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
		.io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
		.io_pmp_1_addr(pmp_io_pmp_1_addr),
		.io_pmp_1_mask(pmp_io_pmp_1_mask),
		.io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
		.io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
		.io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
		.io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
		.io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
		.io_pmp_2_addr(pmp_io_pmp_2_addr),
		.io_pmp_2_mask(pmp_io_pmp_2_mask),
		.io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
		.io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
		.io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
		.io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
		.io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
		.io_pmp_3_addr(pmp_io_pmp_3_addr),
		.io_pmp_3_mask(pmp_io_pmp_3_mask),
		.io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
		.io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
		.io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
		.io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
		.io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
		.io_pmp_4_addr(pmp_io_pmp_4_addr),
		.io_pmp_4_mask(pmp_io_pmp_4_mask),
		.io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
		.io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
		.io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
		.io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
		.io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
		.io_pmp_5_addr(pmp_io_pmp_5_addr),
		.io_pmp_5_mask(pmp_io_pmp_5_mask),
		.io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
		.io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
		.io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
		.io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
		.io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
		.io_pmp_6_addr(pmp_io_pmp_6_addr),
		.io_pmp_6_mask(pmp_io_pmp_6_mask),
		.io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
		.io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
		.io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
		.io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
		.io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
		.io_pmp_7_addr(pmp_io_pmp_7_addr),
		.io_pmp_7_mask(pmp_io_pmp_7_mask),
		.io_addr(pmp_io_addr),
		.io_r(pmp_io_r),
		.io_w(pmp_io_w),
		.io_x(pmp_io_x)
	);
	assign io_resp_paddr = {vpn, io_req_bits_vaddr[11:0]};
	assign io_resp_ae_inst = |_io_resp_ae_inst_T_1;
	assign pmp_io_prv = mpu_priv[1:0];
	assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l;
	assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a;
	assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x;
	assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w;
	assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r;
	assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr;
	assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask;
	assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l;
	assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a;
	assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x;
	assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w;
	assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r;
	assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr;
	assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask;
	assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l;
	assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a;
	assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x;
	assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w;
	assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r;
	assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr;
	assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask;
	assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l;
	assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a;
	assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x;
	assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w;
	assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r;
	assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr;
	assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask;
	assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l;
	assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a;
	assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x;
	assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w;
	assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r;
	assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr;
	assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask;
	assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l;
	assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a;
	assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x;
	assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w;
	assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r;
	assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr;
	assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask;
	assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l;
	assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a;
	assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x;
	assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w;
	assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r;
	assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr;
	assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask;
	assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l;
	assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a;
	assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x;
	assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w;
	assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r;
	assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr;
	assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask;
	assign pmp_io_addr = {mpu_ppn, io_req_bits_vaddr[11:0]};
endmodule
module Frontend (
	clock,
	reset,
	auto_icache_master_out_a_ready,
	auto_icache_master_out_a_valid,
	auto_icache_master_out_a_bits_address,
	auto_icache_master_out_d_valid,
	auto_icache_master_out_d_bits_opcode,
	auto_icache_master_out_d_bits_size,
	auto_icache_master_out_d_bits_data,
	auto_icache_master_out_d_bits_corrupt,
	io_cpu_might_request,
	io_cpu_req_valid,
	io_cpu_req_bits_pc,
	io_cpu_req_bits_speculative,
	io_cpu_resp_ready,
	io_cpu_resp_valid,
	io_cpu_resp_bits_pc,
	io_cpu_resp_bits_data,
	io_cpu_resp_bits_xcpt_ae_inst,
	io_cpu_resp_bits_replay,
	io_cpu_btb_update_valid,
	io_cpu_bht_update_valid,
	io_cpu_flush_icache,
	io_cpu_npc,
	io_ptw_status_debug,
	io_ptw_pmp_0_cfg_l,
	io_ptw_pmp_0_cfg_a,
	io_ptw_pmp_0_cfg_x,
	io_ptw_pmp_0_cfg_w,
	io_ptw_pmp_0_cfg_r,
	io_ptw_pmp_0_addr,
	io_ptw_pmp_0_mask,
	io_ptw_pmp_1_cfg_l,
	io_ptw_pmp_1_cfg_a,
	io_ptw_pmp_1_cfg_x,
	io_ptw_pmp_1_cfg_w,
	io_ptw_pmp_1_cfg_r,
	io_ptw_pmp_1_addr,
	io_ptw_pmp_1_mask,
	io_ptw_pmp_2_cfg_l,
	io_ptw_pmp_2_cfg_a,
	io_ptw_pmp_2_cfg_x,
	io_ptw_pmp_2_cfg_w,
	io_ptw_pmp_2_cfg_r,
	io_ptw_pmp_2_addr,
	io_ptw_pmp_2_mask,
	io_ptw_pmp_3_cfg_l,
	io_ptw_pmp_3_cfg_a,
	io_ptw_pmp_3_cfg_x,
	io_ptw_pmp_3_cfg_w,
	io_ptw_pmp_3_cfg_r,
	io_ptw_pmp_3_addr,
	io_ptw_pmp_3_mask,
	io_ptw_pmp_4_cfg_l,
	io_ptw_pmp_4_cfg_a,
	io_ptw_pmp_4_cfg_x,
	io_ptw_pmp_4_cfg_w,
	io_ptw_pmp_4_cfg_r,
	io_ptw_pmp_4_addr,
	io_ptw_pmp_4_mask,
	io_ptw_pmp_5_cfg_l,
	io_ptw_pmp_5_cfg_a,
	io_ptw_pmp_5_cfg_x,
	io_ptw_pmp_5_cfg_w,
	io_ptw_pmp_5_cfg_r,
	io_ptw_pmp_5_addr,
	io_ptw_pmp_5_mask,
	io_ptw_pmp_6_cfg_l,
	io_ptw_pmp_6_cfg_a,
	io_ptw_pmp_6_cfg_x,
	io_ptw_pmp_6_cfg_w,
	io_ptw_pmp_6_cfg_r,
	io_ptw_pmp_6_addr,
	io_ptw_pmp_6_mask,
	io_ptw_pmp_7_cfg_l,
	io_ptw_pmp_7_cfg_a,
	io_ptw_pmp_7_cfg_x,
	io_ptw_pmp_7_cfg_w,
	io_ptw_pmp_7_cfg_r,
	io_ptw_pmp_7_addr,
	io_ptw_pmp_7_mask,
	io_ptw_customCSRs_csrs_0_value
);
	input clock;
	input reset;
	input auto_icache_master_out_a_ready;
	output wire auto_icache_master_out_a_valid;
	output wire [31:0] auto_icache_master_out_a_bits_address;
	input auto_icache_master_out_d_valid;
	input [2:0] auto_icache_master_out_d_bits_opcode;
	input [3:0] auto_icache_master_out_d_bits_size;
	input [31:0] auto_icache_master_out_d_bits_data;
	input auto_icache_master_out_d_bits_corrupt;
	input io_cpu_might_request;
	input io_cpu_req_valid;
	input [31:0] io_cpu_req_bits_pc;
	input io_cpu_req_bits_speculative;
	input io_cpu_resp_ready;
	output wire io_cpu_resp_valid;
	output wire [31:0] io_cpu_resp_bits_pc;
	output wire [31:0] io_cpu_resp_bits_data;
	output wire io_cpu_resp_bits_xcpt_ae_inst;
	output wire io_cpu_resp_bits_replay;
	input io_cpu_btb_update_valid;
	input io_cpu_bht_update_valid;
	input io_cpu_flush_icache;
	output wire [31:0] io_cpu_npc;
	input io_ptw_status_debug;
	input io_ptw_pmp_0_cfg_l;
	input [1:0] io_ptw_pmp_0_cfg_a;
	input io_ptw_pmp_0_cfg_x;
	input io_ptw_pmp_0_cfg_w;
	input io_ptw_pmp_0_cfg_r;
	input [29:0] io_ptw_pmp_0_addr;
	input [31:0] io_ptw_pmp_0_mask;
	input io_ptw_pmp_1_cfg_l;
	input [1:0] io_ptw_pmp_1_cfg_a;
	input io_ptw_pmp_1_cfg_x;
	input io_ptw_pmp_1_cfg_w;
	input io_ptw_pmp_1_cfg_r;
	input [29:0] io_ptw_pmp_1_addr;
	input [31:0] io_ptw_pmp_1_mask;
	input io_ptw_pmp_2_cfg_l;
	input [1:0] io_ptw_pmp_2_cfg_a;
	input io_ptw_pmp_2_cfg_x;
	input io_ptw_pmp_2_cfg_w;
	input io_ptw_pmp_2_cfg_r;
	input [29:0] io_ptw_pmp_2_addr;
	input [31:0] io_ptw_pmp_2_mask;
	input io_ptw_pmp_3_cfg_l;
	input [1:0] io_ptw_pmp_3_cfg_a;
	input io_ptw_pmp_3_cfg_x;
	input io_ptw_pmp_3_cfg_w;
	input io_ptw_pmp_3_cfg_r;
	input [29:0] io_ptw_pmp_3_addr;
	input [31:0] io_ptw_pmp_3_mask;
	input io_ptw_pmp_4_cfg_l;
	input [1:0] io_ptw_pmp_4_cfg_a;
	input io_ptw_pmp_4_cfg_x;
	input io_ptw_pmp_4_cfg_w;
	input io_ptw_pmp_4_cfg_r;
	input [29:0] io_ptw_pmp_4_addr;
	input [31:0] io_ptw_pmp_4_mask;
	input io_ptw_pmp_5_cfg_l;
	input [1:0] io_ptw_pmp_5_cfg_a;
	input io_ptw_pmp_5_cfg_x;
	input io_ptw_pmp_5_cfg_w;
	input io_ptw_pmp_5_cfg_r;
	input [29:0] io_ptw_pmp_5_addr;
	input [31:0] io_ptw_pmp_5_mask;
	input io_ptw_pmp_6_cfg_l;
	input [1:0] io_ptw_pmp_6_cfg_a;
	input io_ptw_pmp_6_cfg_x;
	input io_ptw_pmp_6_cfg_w;
	input io_ptw_pmp_6_cfg_r;
	input [29:0] io_ptw_pmp_6_addr;
	input [31:0] io_ptw_pmp_6_mask;
	input io_ptw_pmp_7_cfg_l;
	input [1:0] io_ptw_pmp_7_cfg_a;
	input io_ptw_pmp_7_cfg_x;
	input io_ptw_pmp_7_cfg_w;
	input io_ptw_pmp_7_cfg_r;
	input [29:0] io_ptw_pmp_7_addr;
	input [31:0] io_ptw_pmp_7_mask;
	input [31:0] io_ptw_customCSRs_csrs_0_value;
	wire icache_clock;
	wire icache_reset;
	wire icache_auto_master_out_a_ready;
	wire icache_auto_master_out_a_valid;
	wire [31:0] icache_auto_master_out_a_bits_address;
	wire icache_auto_master_out_d_valid;
	wire [2:0] icache_auto_master_out_d_bits_opcode;
	wire [3:0] icache_auto_master_out_d_bits_size;
	wire [31:0] icache_auto_master_out_d_bits_data;
	wire icache_auto_master_out_d_bits_corrupt;
	wire icache_io_req_ready;
	wire icache_io_req_valid;
	wire [31:0] icache_io_req_bits_addr;
	wire [31:0] icache_io_s1_paddr;
	wire icache_io_s1_kill;
	wire icache_io_s2_kill;
	wire icache_io_resp_valid;
	wire [31:0] icache_io_resp_bits_data;
	wire icache_io_resp_bits_ae;
	wire icache_io_invalidate;
	wire fq_clock;
	wire fq_reset;
	wire fq_io_enq_ready;
	wire fq_io_enq_valid;
	wire [31:0] fq_io_enq_bits_pc;
	wire [31:0] fq_io_enq_bits_data;
	wire fq_io_enq_bits_xcpt_ae_inst;
	wire fq_io_enq_bits_replay;
	wire fq_io_deq_ready;
	wire fq_io_deq_valid;
	wire [31:0] fq_io_deq_bits_pc;
	wire [31:0] fq_io_deq_bits_data;
	wire fq_io_deq_bits_xcpt_ae_inst;
	wire fq_io_deq_bits_replay;
	wire [4:0] fq_io_mask;
	wire [31:0] tlb_io_req_bits_vaddr;
	wire [31:0] tlb_io_resp_paddr;
	wire tlb_io_resp_ae_inst;
	wire tlb_io_ptw_status_debug;
	wire tlb_io_ptw_pmp_0_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_0_cfg_a;
	wire tlb_io_ptw_pmp_0_cfg_x;
	wire tlb_io_ptw_pmp_0_cfg_w;
	wire tlb_io_ptw_pmp_0_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_0_addr;
	wire [31:0] tlb_io_ptw_pmp_0_mask;
	wire tlb_io_ptw_pmp_1_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_1_cfg_a;
	wire tlb_io_ptw_pmp_1_cfg_x;
	wire tlb_io_ptw_pmp_1_cfg_w;
	wire tlb_io_ptw_pmp_1_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_1_addr;
	wire [31:0] tlb_io_ptw_pmp_1_mask;
	wire tlb_io_ptw_pmp_2_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_2_cfg_a;
	wire tlb_io_ptw_pmp_2_cfg_x;
	wire tlb_io_ptw_pmp_2_cfg_w;
	wire tlb_io_ptw_pmp_2_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_2_addr;
	wire [31:0] tlb_io_ptw_pmp_2_mask;
	wire tlb_io_ptw_pmp_3_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_3_cfg_a;
	wire tlb_io_ptw_pmp_3_cfg_x;
	wire tlb_io_ptw_pmp_3_cfg_w;
	wire tlb_io_ptw_pmp_3_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_3_addr;
	wire [31:0] tlb_io_ptw_pmp_3_mask;
	wire tlb_io_ptw_pmp_4_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_4_cfg_a;
	wire tlb_io_ptw_pmp_4_cfg_x;
	wire tlb_io_ptw_pmp_4_cfg_w;
	wire tlb_io_ptw_pmp_4_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_4_addr;
	wire [31:0] tlb_io_ptw_pmp_4_mask;
	wire tlb_io_ptw_pmp_5_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_5_cfg_a;
	wire tlb_io_ptw_pmp_5_cfg_x;
	wire tlb_io_ptw_pmp_5_cfg_w;
	wire tlb_io_ptw_pmp_5_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_5_addr;
	wire [31:0] tlb_io_ptw_pmp_5_mask;
	wire tlb_io_ptw_pmp_6_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_6_cfg_a;
	wire tlb_io_ptw_pmp_6_cfg_x;
	wire tlb_io_ptw_pmp_6_cfg_w;
	wire tlb_io_ptw_pmp_6_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_6_addr;
	wire [31:0] tlb_io_ptw_pmp_6_mask;
	wire tlb_io_ptw_pmp_7_cfg_l;
	wire [1:0] tlb_io_ptw_pmp_7_cfg_a;
	wire tlb_io_ptw_pmp_7_cfg_x;
	wire tlb_io_ptw_pmp_7_cfg_w;
	wire tlb_io_ptw_pmp_7_cfg_r;
	wire [29:0] tlb_io_ptw_pmp_7_addr;
	wire [31:0] tlb_io_ptw_pmp_7_mask;
	wire _T_9 = ~reset;
	reg s1_valid;
	reg s2_valid;
	wire _s0_fq_has_space_T_4 = ~s1_valid;
	wire _s0_fq_has_space_T_5 = ~s2_valid;
	wire _s0_fq_has_space_T_7 = ~fq_io_mask[3] & (~s1_valid | ~s2_valid);
	wire _s0_fq_has_space_T_8 = ~fq_io_mask[2] | _s0_fq_has_space_T_7;
	wire _s0_fq_has_space_T_14 = ~fq_io_mask[4] & (_s0_fq_has_space_T_4 & _s0_fq_has_space_T_5);
	wire s0_fq_has_space = _s0_fq_has_space_T_8 | _s0_fq_has_space_T_14;
	wire s0_valid = io_cpu_req_valid | s0_fq_has_space;
	reg [31:0] s1_pc;
	reg s1_speculative;
	reg [31:0] s2_pc;
	reg s2_tlb_resp_ae_inst;
	reg s2_speculative;
	wire [31:0] _s1_base_pc_T = ~s1_pc;
	wire [31:0] _s1_base_pc_T_1 = _s1_base_pc_T | 32'h00000003;
	wire [31:0] s1_base_pc = ~_s1_base_pc_T_1;
	wire [31:0] ntpc = s1_base_pc + 32'h00000004;
	wire _s2_replay_T = fq_io_enq_ready & fq_io_enq_valid;
	reg s2_replay_REG;
	wire s2_replay = (s2_valid & ~_s2_replay_T) | s2_replay_REG;
	wire [31:0] npc = (s2_replay ? s2_pc : ntpc);
	wire s0_speculative = s1_speculative | (s2_valid & ~s2_speculative);
	wire _GEN_0 = ~s2_replay & ~io_cpu_req_valid;
	reg fq_io_enq_valid_REG;
	wire [31:0] _io_cpu_npc_T = (io_cpu_req_valid ? io_cpu_req_bits_pc : npc);
	wire [31:0] _io_cpu_npc_T_1 = ~_io_cpu_npc_T;
	wire [31:0] _io_cpu_npc_T_2 = _io_cpu_npc_T_1 | 32'h00000001;
	ICache icache(
		.clock(icache_clock),
		.reset(icache_reset),
		.auto_master_out_a_ready(icache_auto_master_out_a_ready),
		.auto_master_out_a_valid(icache_auto_master_out_a_valid),
		.auto_master_out_a_bits_address(icache_auto_master_out_a_bits_address),
		.auto_master_out_d_valid(icache_auto_master_out_d_valid),
		.auto_master_out_d_bits_opcode(icache_auto_master_out_d_bits_opcode),
		.auto_master_out_d_bits_size(icache_auto_master_out_d_bits_size),
		.auto_master_out_d_bits_data(icache_auto_master_out_d_bits_data),
		.auto_master_out_d_bits_corrupt(icache_auto_master_out_d_bits_corrupt),
		.io_req_ready(icache_io_req_ready),
		.io_req_valid(icache_io_req_valid),
		.io_req_bits_addr(icache_io_req_bits_addr),
		.io_s1_paddr(icache_io_s1_paddr),
		.io_s1_kill(icache_io_s1_kill),
		.io_s2_kill(icache_io_s2_kill),
		.io_resp_valid(icache_io_resp_valid),
		.io_resp_bits_data(icache_io_resp_bits_data),
		.io_resp_bits_ae(icache_io_resp_bits_ae),
		.io_invalidate(icache_io_invalidate)
	);
	ShiftQueue fq(
		.clock(fq_clock),
		.reset(fq_reset),
		.io_enq_ready(fq_io_enq_ready),
		.io_enq_valid(fq_io_enq_valid),
		.io_enq_bits_pc(fq_io_enq_bits_pc),
		.io_enq_bits_data(fq_io_enq_bits_data),
		.io_enq_bits_xcpt_ae_inst(fq_io_enq_bits_xcpt_ae_inst),
		.io_enq_bits_replay(fq_io_enq_bits_replay),
		.io_deq_ready(fq_io_deq_ready),
		.io_deq_valid(fq_io_deq_valid),
		.io_deq_bits_pc(fq_io_deq_bits_pc),
		.io_deq_bits_data(fq_io_deq_bits_data),
		.io_deq_bits_xcpt_ae_inst(fq_io_deq_bits_xcpt_ae_inst),
		.io_deq_bits_replay(fq_io_deq_bits_replay),
		.io_mask(fq_io_mask)
	);
	TLB_1 tlb(
		.io_req_bits_vaddr(tlb_io_req_bits_vaddr),
		.io_resp_paddr(tlb_io_resp_paddr),
		.io_resp_ae_inst(tlb_io_resp_ae_inst),
		.io_ptw_status_debug(tlb_io_ptw_status_debug),
		.io_ptw_pmp_0_cfg_l(tlb_io_ptw_pmp_0_cfg_l),
		.io_ptw_pmp_0_cfg_a(tlb_io_ptw_pmp_0_cfg_a),
		.io_ptw_pmp_0_cfg_x(tlb_io_ptw_pmp_0_cfg_x),
		.io_ptw_pmp_0_cfg_w(tlb_io_ptw_pmp_0_cfg_w),
		.io_ptw_pmp_0_cfg_r(tlb_io_ptw_pmp_0_cfg_r),
		.io_ptw_pmp_0_addr(tlb_io_ptw_pmp_0_addr),
		.io_ptw_pmp_0_mask(tlb_io_ptw_pmp_0_mask),
		.io_ptw_pmp_1_cfg_l(tlb_io_ptw_pmp_1_cfg_l),
		.io_ptw_pmp_1_cfg_a(tlb_io_ptw_pmp_1_cfg_a),
		.io_ptw_pmp_1_cfg_x(tlb_io_ptw_pmp_1_cfg_x),
		.io_ptw_pmp_1_cfg_w(tlb_io_ptw_pmp_1_cfg_w),
		.io_ptw_pmp_1_cfg_r(tlb_io_ptw_pmp_1_cfg_r),
		.io_ptw_pmp_1_addr(tlb_io_ptw_pmp_1_addr),
		.io_ptw_pmp_1_mask(tlb_io_ptw_pmp_1_mask),
		.io_ptw_pmp_2_cfg_l(tlb_io_ptw_pmp_2_cfg_l),
		.io_ptw_pmp_2_cfg_a(tlb_io_ptw_pmp_2_cfg_a),
		.io_ptw_pmp_2_cfg_x(tlb_io_ptw_pmp_2_cfg_x),
		.io_ptw_pmp_2_cfg_w(tlb_io_ptw_pmp_2_cfg_w),
		.io_ptw_pmp_2_cfg_r(tlb_io_ptw_pmp_2_cfg_r),
		.io_ptw_pmp_2_addr(tlb_io_ptw_pmp_2_addr),
		.io_ptw_pmp_2_mask(tlb_io_ptw_pmp_2_mask),
		.io_ptw_pmp_3_cfg_l(tlb_io_ptw_pmp_3_cfg_l),
		.io_ptw_pmp_3_cfg_a(tlb_io_ptw_pmp_3_cfg_a),
		.io_ptw_pmp_3_cfg_x(tlb_io_ptw_pmp_3_cfg_x),
		.io_ptw_pmp_3_cfg_w(tlb_io_ptw_pmp_3_cfg_w),
		.io_ptw_pmp_3_cfg_r(tlb_io_ptw_pmp_3_cfg_r),
		.io_ptw_pmp_3_addr(tlb_io_ptw_pmp_3_addr),
		.io_ptw_pmp_3_mask(tlb_io_ptw_pmp_3_mask),
		.io_ptw_pmp_4_cfg_l(tlb_io_ptw_pmp_4_cfg_l),
		.io_ptw_pmp_4_cfg_a(tlb_io_ptw_pmp_4_cfg_a),
		.io_ptw_pmp_4_cfg_x(tlb_io_ptw_pmp_4_cfg_x),
		.io_ptw_pmp_4_cfg_w(tlb_io_ptw_pmp_4_cfg_w),
		.io_ptw_pmp_4_cfg_r(tlb_io_ptw_pmp_4_cfg_r),
		.io_ptw_pmp_4_addr(tlb_io_ptw_pmp_4_addr),
		.io_ptw_pmp_4_mask(tlb_io_ptw_pmp_4_mask),
		.io_ptw_pmp_5_cfg_l(tlb_io_ptw_pmp_5_cfg_l),
		.io_ptw_pmp_5_cfg_a(tlb_io_ptw_pmp_5_cfg_a),
		.io_ptw_pmp_5_cfg_x(tlb_io_ptw_pmp_5_cfg_x),
		.io_ptw_pmp_5_cfg_w(tlb_io_ptw_pmp_5_cfg_w),
		.io_ptw_pmp_5_cfg_r(tlb_io_ptw_pmp_5_cfg_r),
		.io_ptw_pmp_5_addr(tlb_io_ptw_pmp_5_addr),
		.io_ptw_pmp_5_mask(tlb_io_ptw_pmp_5_mask),
		.io_ptw_pmp_6_cfg_l(tlb_io_ptw_pmp_6_cfg_l),
		.io_ptw_pmp_6_cfg_a(tlb_io_ptw_pmp_6_cfg_a),
		.io_ptw_pmp_6_cfg_x(tlb_io_ptw_pmp_6_cfg_x),
		.io_ptw_pmp_6_cfg_w(tlb_io_ptw_pmp_6_cfg_w),
		.io_ptw_pmp_6_cfg_r(tlb_io_ptw_pmp_6_cfg_r),
		.io_ptw_pmp_6_addr(tlb_io_ptw_pmp_6_addr),
		.io_ptw_pmp_6_mask(tlb_io_ptw_pmp_6_mask),
		.io_ptw_pmp_7_cfg_l(tlb_io_ptw_pmp_7_cfg_l),
		.io_ptw_pmp_7_cfg_a(tlb_io_ptw_pmp_7_cfg_a),
		.io_ptw_pmp_7_cfg_x(tlb_io_ptw_pmp_7_cfg_x),
		.io_ptw_pmp_7_cfg_w(tlb_io_ptw_pmp_7_cfg_w),
		.io_ptw_pmp_7_cfg_r(tlb_io_ptw_pmp_7_cfg_r),
		.io_ptw_pmp_7_addr(tlb_io_ptw_pmp_7_addr),
		.io_ptw_pmp_7_mask(tlb_io_ptw_pmp_7_mask)
	);
	assign auto_icache_master_out_a_valid = icache_auto_master_out_a_valid;
	assign auto_icache_master_out_a_bits_address = icache_auto_master_out_a_bits_address;
	assign io_cpu_resp_valid = fq_io_deq_valid;
	assign io_cpu_resp_bits_pc = fq_io_deq_bits_pc;
	assign io_cpu_resp_bits_data = fq_io_deq_bits_data;
	assign io_cpu_resp_bits_xcpt_ae_inst = fq_io_deq_bits_xcpt_ae_inst;
	assign io_cpu_resp_bits_replay = fq_io_deq_bits_replay;
	assign io_cpu_npc = ~_io_cpu_npc_T_2;
	assign icache_clock = clock;
	assign icache_reset = reset;
	assign icache_auto_master_out_a_ready = auto_icache_master_out_a_ready;
	assign icache_auto_master_out_d_valid = auto_icache_master_out_d_valid;
	assign icache_auto_master_out_d_bits_opcode = auto_icache_master_out_d_bits_opcode;
	assign icache_auto_master_out_d_bits_size = auto_icache_master_out_d_bits_size;
	assign icache_auto_master_out_d_bits_data = auto_icache_master_out_d_bits_data;
	assign icache_auto_master_out_d_bits_corrupt = auto_icache_master_out_d_bits_corrupt;
	assign icache_io_req_valid = io_cpu_req_valid | s0_fq_has_space;
	assign icache_io_req_bits_addr = io_cpu_npc;
	assign icache_io_s1_paddr = tlb_io_resp_paddr;
	assign icache_io_s1_kill = io_cpu_req_valid | s2_replay;
	assign icache_io_s2_kill = s2_speculative | s2_tlb_resp_ae_inst;
	assign icache_io_invalidate = io_cpu_flush_icache;
	assign fq_clock = clock;
	assign fq_reset = reset | io_cpu_req_valid;
	assign fq_io_enq_valid = (fq_io_enq_valid_REG & s2_valid) & (icache_io_resp_valid | icache_io_s2_kill);
	assign fq_io_enq_bits_pc = s2_pc;
	assign fq_io_enq_bits_data = icache_io_resp_bits_data;
	assign fq_io_enq_bits_xcpt_ae_inst = (icache_io_resp_valid & icache_io_resp_bits_ae) | s2_tlb_resp_ae_inst;
	assign fq_io_enq_bits_replay = (icache_io_s2_kill & ~icache_io_resp_valid) & ~s2_tlb_resp_ae_inst;
	assign fq_io_deq_ready = io_cpu_resp_ready;
	assign tlb_io_req_bits_vaddr = s1_pc;
	assign tlb_io_ptw_status_debug = io_ptw_status_debug;
	assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l;
	assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a;
	assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x;
	assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w;
	assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r;
	assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr;
	assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask;
	assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l;
	assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a;
	assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x;
	assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w;
	assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r;
	assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr;
	assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask;
	assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l;
	assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a;
	assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x;
	assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w;
	assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r;
	assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr;
	assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask;
	assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l;
	assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a;
	assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x;
	assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w;
	assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r;
	assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr;
	assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask;
	assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l;
	assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a;
	assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x;
	assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w;
	assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r;
	assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr;
	assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask;
	assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l;
	assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a;
	assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x;
	assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w;
	assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r;
	assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr;
	assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask;
	assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l;
	assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a;
	assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x;
	assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w;
	assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r;
	assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr;
	assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask;
	assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l;
	assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a;
	assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x;
	assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w;
	assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r;
	assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr;
	assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask;
	always @(posedge clock) begin
		s1_valid <= io_cpu_req_valid | s0_fq_has_space;
		if (reset)
			s2_valid <= 1'h0;
		else
			s2_valid <= _GEN_0;
		s1_pc <= io_cpu_npc;
		if (io_cpu_req_valid)
			s1_speculative <= io_cpu_req_bits_speculative;
		else if (s2_replay)
			s1_speculative <= s2_speculative;
		else
			s1_speculative <= s0_speculative;
		if (reset)
			s2_pc <= 32'h00010040;
		else if (~s2_replay)
			s2_pc <= s1_pc;
		if (~s2_replay)
			s2_tlb_resp_ae_inst <= tlb_io_resp_ae_inst;
		if (reset)
			s2_speculative <= 1'h0;
		else if (~s2_replay)
			s2_speculative <= s1_speculative;
		s2_replay_REG <= reset | (s2_replay & ~s0_valid);
		fq_io_enq_valid_REG <= s1_valid;
	end
endmodule
module ScratchpadSlavePort (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	io_dmem_req_ready,
	io_dmem_req_valid,
	io_dmem_req_bits_addr,
	io_dmem_req_bits_cmd,
	io_dmem_req_bits_size,
	io_dmem_s1_kill,
	io_dmem_s1_data_data,
	io_dmem_s1_data_mask,
	io_dmem_s2_nack,
	io_dmem_resp_valid,
	io_dmem_resp_bits_data_raw
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [1:0] auto_in_a_bits_size;
	input [8:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_size;
	output wire [8:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input io_dmem_req_ready;
	output wire io_dmem_req_valid;
	output wire [31:0] io_dmem_req_bits_addr;
	output wire [4:0] io_dmem_req_bits_cmd;
	output wire [1:0] io_dmem_req_bits_size;
	output wire io_dmem_s1_kill;
	output wire [31:0] io_dmem_s1_data_data;
	output wire [3:0] io_dmem_s1_data_mask;
	input io_dmem_s2_nack;
	input io_dmem_resp_valid;
	input [31:0] io_dmem_resp_bits_data_raw;
	reg [2:0] state;
	wire [2:0] _GEN_0 = (state == 3'h1 ? 3'h2 : state);
	wire _T_1 = state == 3'h4;
	wire [2:0] _GEN_1 = ((state == 3'h4) & auto_in_a_valid ? 3'h0 : _GEN_0);
	wire [2:0] _GEN_2 = (io_dmem_resp_valid ? 3'h5 : _GEN_1);
	wire tl_in_d_valid = io_dmem_resp_valid | (state == 3'h5);
	wire _T_3 = auto_in_d_ready & tl_in_d_valid;
	wire _ready_T = state == 3'h0;
	wire _ready_T_1 = state == 3'h2;
	wire ready = (state == 3'h0) | (((state == 3'h2) & io_dmem_resp_valid) & auto_in_d_ready);
	wire _dmem_req_valid_T_1 = state == 3'h3;
	wire dmem_req_valid = (auto_in_a_valid & ready) | (state == 3'h3);
	reg [2:0] acq_opcode;
	reg [2:0] acq_param;
	reg [1:0] acq_size;
	reg [8:0] acq_source;
	reg [31:0] acq_address;
	reg [3:0] acq_mask;
	reg [31:0] acq_data;
	wire tl_in_a_ready = io_dmem_req_ready & ready;
	wire _T_5 = tl_in_a_ready & auto_in_a_valid;
	wire ready_likely = _ready_T | _ready_T_1;
	wire [2:0] _io_dmem_req_bits_T_1_opcode = (_dmem_req_valid_T_1 ? acq_opcode : auto_in_a_bits_opcode);
	wire [2:0] _io_dmem_req_bits_T_1_param = (_dmem_req_valid_T_1 ? acq_param : auto_in_a_bits_param);
	wire [1:0] io_dmem_req_bits_mask_full_desired_mask_size = (_dmem_req_valid_T_1 ? acq_size : auto_in_a_bits_size);
	wire [31:0] io_dmem_req_bits_req_addr = (_dmem_req_valid_T_1 ? acq_address : auto_in_a_bits_address);
	wire [3:0] _io_dmem_req_bits_T_1_mask = (_dmem_req_valid_T_1 ? acq_mask : auto_in_a_bits_mask);
	wire [3:0] _io_dmem_req_bits_req_cmd_T_1 = (3'h0 == _io_dmem_req_bits_T_1_param ? 4'hc : 4'h0);
	wire [3:0] _io_dmem_req_bits_req_cmd_T_3 = (3'h1 == _io_dmem_req_bits_T_1_param ? 4'hd : _io_dmem_req_bits_req_cmd_T_1);
	wire [3:0] _io_dmem_req_bits_req_cmd_T_5 = (3'h2 == _io_dmem_req_bits_T_1_param ? 4'he : _io_dmem_req_bits_req_cmd_T_3);
	wire [3:0] _io_dmem_req_bits_req_cmd_T_7 = (3'h3 == _io_dmem_req_bits_T_1_param ? 4'hf : _io_dmem_req_bits_req_cmd_T_5);
	wire [3:0] _io_dmem_req_bits_req_cmd_T_9 = (3'h4 == _io_dmem_req_bits_T_1_param ? 4'h8 : _io_dmem_req_bits_req_cmd_T_7);
	wire [3:0] _io_dmem_req_bits_req_cmd_T_11 = (3'h0 == _io_dmem_req_bits_T_1_param ? 4'h9 : 4'h0);
	wire [3:0] _io_dmem_req_bits_req_cmd_T_13 = (3'h1 == _io_dmem_req_bits_T_1_param ? 4'ha : _io_dmem_req_bits_req_cmd_T_11);
	wire [3:0] _io_dmem_req_bits_req_cmd_T_15 = (3'h2 == _io_dmem_req_bits_T_1_param ? 4'hb : _io_dmem_req_bits_req_cmd_T_13);
	wire [3:0] _io_dmem_req_bits_req_cmd_T_17 = (3'h3 == _io_dmem_req_bits_T_1_param ? 4'h4 : _io_dmem_req_bits_req_cmd_T_15);
	wire [4:0] _io_dmem_req_bits_req_cmd_T_21 = (3'h1 == _io_dmem_req_bits_T_1_opcode ? 5'h11 : {4'd0, 3'h0 == _io_dmem_req_bits_T_1_opcode});
	wire [4:0] _io_dmem_req_bits_req_cmd_T_23 = (3'h2 == _io_dmem_req_bits_T_1_opcode ? {1'd0, _io_dmem_req_bits_req_cmd_T_9} : _io_dmem_req_bits_req_cmd_T_21);
	wire [4:0] _io_dmem_req_bits_req_cmd_T_25 = (3'h3 == _io_dmem_req_bits_T_1_opcode ? {1'd0, _io_dmem_req_bits_req_cmd_T_17} : _io_dmem_req_bits_req_cmd_T_23);
	wire [4:0] _io_dmem_req_bits_req_cmd_T_27 = (3'h4 == _io_dmem_req_bits_T_1_opcode ? 5'h00 : _io_dmem_req_bits_req_cmd_T_25);
	wire io_dmem_req_bits_mask_full_desired_mask_upper = io_dmem_req_bits_req_addr[0] | (io_dmem_req_bits_mask_full_desired_mask_size >= 2'h1);
	wire io_dmem_req_bits_mask_full_desired_mask_lower = (io_dmem_req_bits_req_addr[0] ? 1'h0 : 1'h1);
	wire [1:0] _io_dmem_req_bits_mask_full_desired_mask_T = {io_dmem_req_bits_mask_full_desired_mask_upper, io_dmem_req_bits_mask_full_desired_mask_lower};
	wire [1:0] _io_dmem_req_bits_mask_full_desired_mask_upper_T_5 = (io_dmem_req_bits_req_addr[1] ? _io_dmem_req_bits_mask_full_desired_mask_T : 2'h0);
	wire [1:0] _io_dmem_req_bits_mask_full_desired_mask_upper_T_7 = (io_dmem_req_bits_mask_full_desired_mask_size >= 2'h2 ? 2'h3 : 2'h0);
	wire [1:0] io_dmem_req_bits_mask_full_desired_mask_upper_1 = _io_dmem_req_bits_mask_full_desired_mask_upper_T_5 | _io_dmem_req_bits_mask_full_desired_mask_upper_T_7;
	wire [1:0] io_dmem_req_bits_mask_full_desired_mask_lower_1 = (io_dmem_req_bits_req_addr[1] ? 2'h0 : _io_dmem_req_bits_mask_full_desired_mask_T);
	wire [3:0] io_dmem_req_bits_mask_full_desired_mask = {io_dmem_req_bits_mask_full_desired_mask_upper_1, io_dmem_req_bits_mask_full_desired_mask_lower_1};
	wire [3:0] _io_dmem_req_bits_mask_full_T = ~io_dmem_req_bits_mask_full_desired_mask;
	wire [3:0] _io_dmem_req_bits_mask_full_T_1 = _io_dmem_req_bits_T_1_mask | _io_dmem_req_bits_mask_full_T;
	wire io_dmem_req_bits_mask_full = &_io_dmem_req_bits_mask_full_T_1;
	wire _bundleIn_0_d_bits_T = acq_opcode == 3'h0;
	wire _bundleIn_0_d_bits_T_1 = acq_opcode == 3'h1;
	wire _bundleIn_0_d_bits_T_2 = _bundleIn_0_d_bits_T | _bundleIn_0_d_bits_T_1;
	reg [31:0] bundleIn_0_d_bits_data_r;
	assign auto_in_a_ready = io_dmem_req_ready & ready;
	assign auto_in_d_valid = io_dmem_resp_valid | (state == 3'h5);
	assign auto_in_d_bits_opcode = (_bundleIn_0_d_bits_T_2 ? 3'h0 : 3'h1);
	assign auto_in_d_bits_size = acq_size;
	assign auto_in_d_bits_source = acq_source;
	assign auto_in_d_bits_data = (_ready_T_1 ? io_dmem_resp_bits_data_raw : bundleIn_0_d_bits_data_r);
	assign io_dmem_req_valid = (auto_in_a_valid & ready_likely) | _dmem_req_valid_T_1;
	assign io_dmem_req_bits_addr = (_dmem_req_valid_T_1 ? acq_address : auto_in_a_bits_address);
	assign io_dmem_req_bits_cmd = (_T_1 | ((_io_dmem_req_bits_T_1_opcode == 3'h1) & io_dmem_req_bits_mask_full) ? 5'h01 : _io_dmem_req_bits_req_cmd_T_27);
	assign io_dmem_req_bits_size = (_dmem_req_valid_T_1 ? acq_size : auto_in_a_bits_size);
	assign io_dmem_s1_kill = state != 3'h1;
	assign io_dmem_s1_data_data = acq_data;
	assign io_dmem_s1_data_mask = acq_mask;
	always @(posedge clock) begin
		if (reset)
			state <= 3'h4;
		else if (dmem_req_valid & io_dmem_req_ready)
			state <= 3'h1;
		else if (io_dmem_s2_nack)
			state <= 3'h3;
		else if (_T_3)
			state <= 3'h0;
		else
			state <= _GEN_2;
		if (_T_5)
			acq_opcode <= auto_in_a_bits_opcode;
		if (_T_5)
			acq_param <= auto_in_a_bits_param;
		if (_T_5)
			acq_size <= auto_in_a_bits_size;
		if (_T_5)
			acq_source <= auto_in_a_bits_source;
		if (_T_5)
			acq_address <= auto_in_a_bits_address;
		if (_T_5)
			acq_mask <= auto_in_a_bits_mask;
		if (_T_5)
			acq_data <= auto_in_a_bits_data;
		if (_ready_T_1)
			bundleIn_0_d_bits_data_r <= io_dmem_resp_bits_data_raw;
	end
endmodule
module Repeater_9 (
	clock,
	reset,
	io_repeat,
	io_full,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask
);
	input clock;
	input reset;
	input io_repeat;
	output wire io_full;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [31:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [31:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	reg full;
	reg [2:0] saved_opcode;
	reg [2:0] saved_param;
	reg [2:0] saved_size;
	reg [2:0] saved_source;
	reg [31:0] saved_address;
	reg [3:0] saved_mask;
	wire _T = io_enq_ready & io_enq_valid;
	wire _GEN_0 = (_T & io_repeat) | full;
	wire _T_2 = io_deq_ready & io_deq_valid;
	assign io_full = full;
	assign io_enq_ready = io_deq_ready & ~full;
	assign io_deq_valid = io_enq_valid | full;
	assign io_deq_bits_opcode = (full ? saved_opcode : io_enq_bits_opcode);
	assign io_deq_bits_param = (full ? saved_param : io_enq_bits_param);
	assign io_deq_bits_size = (full ? saved_size : io_enq_bits_size);
	assign io_deq_bits_source = (full ? saved_source : io_enq_bits_source);
	assign io_deq_bits_address = (full ? saved_address : io_enq_bits_address);
	assign io_deq_bits_mask = (full ? saved_mask : io_enq_bits_mask);
	always @(posedge clock) begin
		if (reset)
			full <= 1'h0;
		else if (_T_2 & ~io_repeat)
			full <= 1'h0;
		else
			full <= _GEN_0;
		if (_T & io_repeat)
			saved_opcode <= io_enq_bits_opcode;
		if (_T & io_repeat)
			saved_param <= io_enq_bits_param;
		if (_T & io_repeat)
			saved_size <= io_enq_bits_size;
		if (_T & io_repeat)
			saved_source <= io_enq_bits_source;
		if (_T & io_repeat)
			saved_address <= io_enq_bits_address;
		if (_T & io_repeat)
			saved_mask <= io_enq_bits_mask;
	end
endmodule
module TLFragmenter_9 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire [8:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_size;
	input [8:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	wire repeater_clock;
	wire repeater_reset;
	wire repeater_io_repeat;
	wire repeater_io_full;
	wire repeater_io_enq_ready;
	wire repeater_io_enq_valid;
	wire [2:0] repeater_io_enq_bits_opcode;
	wire [2:0] repeater_io_enq_bits_param;
	wire [2:0] repeater_io_enq_bits_size;
	wire [2:0] repeater_io_enq_bits_source;
	wire [31:0] repeater_io_enq_bits_address;
	wire [3:0] repeater_io_enq_bits_mask;
	wire repeater_io_deq_ready;
	wire repeater_io_deq_valid;
	wire [2:0] repeater_io_deq_bits_opcode;
	wire [2:0] repeater_io_deq_bits_param;
	wire [2:0] repeater_io_deq_bits_size;
	wire [2:0] repeater_io_deq_bits_source;
	wire [31:0] repeater_io_deq_bits_address;
	wire [3:0] repeater_io_deq_bits_mask;
	reg [3:0] acknum;
	reg [2:0] dOrig;
	reg dToggle;
	wire [3:0] dFragnum = auto_out_d_bits_source[3:0];
	wire dFirst = acknum == 4'h0;
	wire dLast = dFragnum == 4'h0;
	wire [3:0] _dsizeOH_T = 4'h1 << auto_out_d_bits_size;
	wire [2:0] dsizeOH = _dsizeOH_T[2:0];
	wire [4:0] _dsizeOH1_T_1 = 5'h03 << auto_out_d_bits_size;
	wire [1:0] dsizeOH1 = ~_dsizeOH1_T_1[1:0];
	wire dHasData = auto_out_d_bits_opcode[0];
	wire _T_5 = ~reset;
	wire ack_decrement = dHasData | dsizeOH[2];
	wire [5:0] _dFirst_size_T = {dFragnum, 2'h0};
	wire [5:0] _GEN_7 = {4'd0, dsizeOH1};
	wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7;
	wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0};
	wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h01;
	wire [6:0] _dFirst_size_T_4 = {1'h0, _dFirst_size_T_1};
	wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4;
	wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5;
	wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4];
	wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0];
	wire _dFirst_size_T_7 = |dFirst_size_hi;
	wire [3:0] _GEN_8 = {1'd0, dFirst_size_hi};
	wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo;
	wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2];
	wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0];
	wire _dFirst_size_T_9 = |dFirst_size_hi_1;
	wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1;
	wire [2:0] dFirst_size = {_dFirst_size_T_7, _dFirst_size_T_9, _dFirst_size_T_10[1]};
	wire doEarlyAck = auto_out_d_bits_source[5];
	wire _drop_T_1 = (doEarlyAck ? dFirst : dLast);
	wire drop = ~dHasData & ~_drop_T_1;
	wire bundleOut_0_d_ready = auto_in_d_ready | drop;
	wire _T_7 = bundleOut_0_d_ready & auto_out_d_valid;
	wire [3:0] _GEN_9 = {3'd0, ack_decrement};
	wire [3:0] _acknum_T_1 = acknum - _GEN_9;
	wire [2:0] aFrag = (repeater_io_deq_bits_size > 3'h2 ? 3'h2 : repeater_io_deq_bits_size);
	wire [12:0] _aOrigOH1_T_1 = 13'h003f << repeater_io_deq_bits_size;
	wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0];
	wire [8:0] _aFragOH1_T_1 = 9'h003 << aFrag;
	wire [1:0] aFragOH1 = ~_aFragOH1_T_1[1:0];
	wire aHasData = ~repeater_io_deq_bits_opcode[2];
	reg [3:0] gennum;
	wire aFirst = gennum == 4'h0;
	wire [3:0] _old_gennum1_T_2 = gennum - 4'h1;
	wire [3:0] old_gennum1 = (aFirst ? aOrigOH1[5:2] : _old_gennum1_T_2);
	wire [3:0] _new_gennum_T = ~old_gennum1;
	wire [3:0] new_gennum = ~_new_gennum_T;
	reg aToggle_r;
	wire _GEN_5 = (aFirst ? dToggle : aToggle_r);
	wire aToggle = ~_GEN_5;
	wire aFull = repeater_io_deq_bits_opcode == 3'h0;
	wire bundleOut_0_a_valid = repeater_io_deq_valid;
	wire _T_8 = auto_out_a_ready & bundleOut_0_a_valid;
	wire _repeater_io_repeat_T = ~aHasData;
	wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 2'h0};
	wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1;
	wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1;
	wire [5:0] _GEN_10 = {4'd0, aFragOH1};
	wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10;
	wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h03;
	wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4;
	wire [31:0] _GEN_11 = {26'd0, _bundleOut_0_a_bits_address_T_5};
	wire [4:0] bundleOut_0_a_bits_source_lo = {aToggle, new_gennum};
	wire [3:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source, aFull};
	wire _T_9 = ~repeater_io_full;
	Repeater_9 repeater(
		.clock(repeater_clock),
		.reset(repeater_reset),
		.io_repeat(repeater_io_repeat),
		.io_full(repeater_io_full),
		.io_enq_ready(repeater_io_enq_ready),
		.io_enq_valid(repeater_io_enq_valid),
		.io_enq_bits_opcode(repeater_io_enq_bits_opcode),
		.io_enq_bits_param(repeater_io_enq_bits_param),
		.io_enq_bits_size(repeater_io_enq_bits_size),
		.io_enq_bits_source(repeater_io_enq_bits_source),
		.io_enq_bits_address(repeater_io_enq_bits_address),
		.io_enq_bits_mask(repeater_io_enq_bits_mask),
		.io_deq_ready(repeater_io_deq_ready),
		.io_deq_valid(repeater_io_deq_valid),
		.io_deq_bits_opcode(repeater_io_deq_bits_opcode),
		.io_deq_bits_param(repeater_io_deq_bits_param),
		.io_deq_bits_size(repeater_io_deq_bits_size),
		.io_deq_bits_source(repeater_io_deq_bits_source),
		.io_deq_bits_address(repeater_io_deq_bits_address),
		.io_deq_bits_mask(repeater_io_deq_bits_mask)
	);
	assign auto_in_a_ready = repeater_io_enq_ready;
	assign auto_in_d_valid = auto_out_d_valid & ~drop;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_size = (dFirst ? dFirst_size : dOrig);
	assign auto_in_d_bits_source = auto_out_d_bits_source[8:6];
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_out_a_valid = repeater_io_deq_valid;
	assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode;
	assign auto_out_a_bits_param = repeater_io_deq_bits_param;
	assign auto_out_a_bits_size = aFrag[1:0];
	assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi, bundleOut_0_a_bits_source_lo};
	assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11;
	assign auto_out_a_bits_mask = (repeater_io_full ? 4'hf : auto_in_a_bits_mask);
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_d_ready = auto_in_d_ready | drop;
	assign repeater_clock = clock;
	assign repeater_reset = reset;
	assign repeater_io_repeat = ~aHasData & (new_gennum != 4'h0);
	assign repeater_io_enq_valid = auto_in_a_valid;
	assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign repeater_io_enq_bits_param = auto_in_a_bits_param;
	assign repeater_io_enq_bits_size = auto_in_a_bits_size;
	assign repeater_io_enq_bits_source = auto_in_a_bits_source;
	assign repeater_io_enq_bits_address = auto_in_a_bits_address;
	assign repeater_io_enq_bits_mask = auto_in_a_bits_mask;
	assign repeater_io_deq_ready = auto_out_a_ready;
	always @(posedge clock) begin
		if (reset)
			acknum <= 4'h0;
		else if (_T_7)
			if (dFirst)
				acknum <= dFragnum;
			else
				acknum <= _acknum_T_1;
		if (_T_7)
			if (dFirst)
				dOrig <= dFirst_size;
		if (reset)
			dToggle <= 1'h0;
		else if (_T_7)
			if (dFirst)
				dToggle <= auto_out_d_bits_source[4];
		if (reset)
			gennum <= 4'h0;
		else if (_T_8)
			gennum <= new_gennum;
		if (aFirst)
			aToggle_r <= dToggle;
	end
endmodule
module HellaCacheArbiter (
	clock,
	io_requestor_0_req_ready,
	io_requestor_0_req_valid,
	io_requestor_0_req_bits_addr,
	io_requestor_0_req_bits_tag,
	io_requestor_0_req_bits_cmd,
	io_requestor_0_req_bits_size,
	io_requestor_0_req_bits_signed,
	io_requestor_0_s1_kill,
	io_requestor_0_s1_data_data,
	io_requestor_0_s2_nack,
	io_requestor_0_resp_valid,
	io_requestor_0_resp_bits_tag,
	io_requestor_0_resp_bits_data,
	io_requestor_0_resp_bits_replay,
	io_requestor_0_resp_bits_has_data,
	io_requestor_0_resp_bits_data_word_bypass,
	io_requestor_0_replay_next,
	io_requestor_0_s2_xcpt_ma_ld,
	io_requestor_0_s2_xcpt_ma_st,
	io_requestor_0_s2_xcpt_pf_ld,
	io_requestor_0_s2_xcpt_pf_st,
	io_requestor_0_s2_xcpt_ae_ld,
	io_requestor_0_s2_xcpt_ae_st,
	io_requestor_0_ordered,
	io_requestor_0_perf_grant,
	io_requestor_1_req_ready,
	io_requestor_1_req_valid,
	io_requestor_1_req_bits_addr,
	io_requestor_1_req_bits_cmd,
	io_requestor_1_req_bits_size,
	io_requestor_1_s1_kill,
	io_requestor_1_s1_data_data,
	io_requestor_1_s1_data_mask,
	io_requestor_1_s2_nack,
	io_requestor_1_resp_valid,
	io_requestor_1_resp_bits_data_raw,
	io_mem_req_ready,
	io_mem_req_valid,
	io_mem_req_bits_addr,
	io_mem_req_bits_tag,
	io_mem_req_bits_cmd,
	io_mem_req_bits_size,
	io_mem_req_bits_signed,
	io_mem_req_bits_dprv,
	io_mem_req_bits_no_xcpt,
	io_mem_s1_kill,
	io_mem_s1_data_data,
	io_mem_s1_data_mask,
	io_mem_s2_nack,
	io_mem_resp_valid,
	io_mem_resp_bits_tag,
	io_mem_resp_bits_data,
	io_mem_resp_bits_replay,
	io_mem_resp_bits_has_data,
	io_mem_resp_bits_data_word_bypass,
	io_mem_resp_bits_data_raw,
	io_mem_replay_next,
	io_mem_s2_xcpt_ma_ld,
	io_mem_s2_xcpt_ma_st,
	io_mem_s2_xcpt_pf_ld,
	io_mem_s2_xcpt_pf_st,
	io_mem_s2_xcpt_ae_ld,
	io_mem_s2_xcpt_ae_st,
	io_mem_ordered,
	io_mem_perf_grant
);
	input clock;
	output wire io_requestor_0_req_ready;
	input io_requestor_0_req_valid;
	input [31:0] io_requestor_0_req_bits_addr;
	input [6:0] io_requestor_0_req_bits_tag;
	input [4:0] io_requestor_0_req_bits_cmd;
	input [1:0] io_requestor_0_req_bits_size;
	input io_requestor_0_req_bits_signed;
	input io_requestor_0_s1_kill;
	input [31:0] io_requestor_0_s1_data_data;
	output wire io_requestor_0_s2_nack;
	output wire io_requestor_0_resp_valid;
	output wire [6:0] io_requestor_0_resp_bits_tag;
	output wire [31:0] io_requestor_0_resp_bits_data;
	output wire io_requestor_0_resp_bits_replay;
	output wire io_requestor_0_resp_bits_has_data;
	output wire [31:0] io_requestor_0_resp_bits_data_word_bypass;
	output wire io_requestor_0_replay_next;
	output wire io_requestor_0_s2_xcpt_ma_ld;
	output wire io_requestor_0_s2_xcpt_ma_st;
	output wire io_requestor_0_s2_xcpt_pf_ld;
	output wire io_requestor_0_s2_xcpt_pf_st;
	output wire io_requestor_0_s2_xcpt_ae_ld;
	output wire io_requestor_0_s2_xcpt_ae_st;
	output wire io_requestor_0_ordered;
	output wire io_requestor_0_perf_grant;
	output wire io_requestor_1_req_ready;
	input io_requestor_1_req_valid;
	input [31:0] io_requestor_1_req_bits_addr;
	input [4:0] io_requestor_1_req_bits_cmd;
	input [1:0] io_requestor_1_req_bits_size;
	input io_requestor_1_s1_kill;
	input [31:0] io_requestor_1_s1_data_data;
	input [3:0] io_requestor_1_s1_data_mask;
	output wire io_requestor_1_s2_nack;
	output wire io_requestor_1_resp_valid;
	output wire [31:0] io_requestor_1_resp_bits_data_raw;
	input io_mem_req_ready;
	output wire io_mem_req_valid;
	output wire [31:0] io_mem_req_bits_addr;
	output wire [6:0] io_mem_req_bits_tag;
	output wire [4:0] io_mem_req_bits_cmd;
	output wire [1:0] io_mem_req_bits_size;
	output wire io_mem_req_bits_signed;
	output wire [1:0] io_mem_req_bits_dprv;
	output wire io_mem_req_bits_no_xcpt;
	output wire io_mem_s1_kill;
	output wire [31:0] io_mem_s1_data_data;
	output wire [3:0] io_mem_s1_data_mask;
	input io_mem_s2_nack;
	input io_mem_resp_valid;
	input [6:0] io_mem_resp_bits_tag;
	input [31:0] io_mem_resp_bits_data;
	input io_mem_resp_bits_replay;
	input io_mem_resp_bits_has_data;
	input [31:0] io_mem_resp_bits_data_word_bypass;
	input [31:0] io_mem_resp_bits_data_raw;
	input io_mem_replay_next;
	input io_mem_s2_xcpt_ma_ld;
	input io_mem_s2_xcpt_ma_st;
	input io_mem_s2_xcpt_pf_ld;
	input io_mem_s2_xcpt_pf_st;
	input io_mem_s2_xcpt_ae_ld;
	input io_mem_s2_xcpt_ae_st;
	input io_mem_ordered;
	input io_mem_perf_grant;
	reg s1_id;
	reg s2_id;
	wire [7:0] _io_mem_req_bits_tag_T_1 = {io_requestor_0_req_bits_tag, 1'h0};
	wire [7:0] _GEN_1 = (io_requestor_0_req_valid ? _io_mem_req_bits_tag_T_1 : 8'h01);
	wire _T_1 = ~s2_id;
	wire tag_hit = ~io_mem_resp_bits_tag[0];
	assign io_requestor_0_req_ready = io_mem_req_ready;
	assign io_requestor_0_s2_nack = io_mem_s2_nack & _T_1;
	assign io_requestor_0_resp_valid = io_mem_resp_valid & tag_hit;
	assign io_requestor_0_resp_bits_tag = {1'd0, io_mem_resp_bits_tag[6:1]};
	assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
	assign io_requestor_0_resp_bits_replay = io_mem_resp_bits_replay;
	assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
	assign io_requestor_0_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
	assign io_requestor_0_replay_next = io_mem_replay_next;
	assign io_requestor_0_s2_xcpt_ma_ld = io_mem_s2_xcpt_ma_ld;
	assign io_requestor_0_s2_xcpt_ma_st = io_mem_s2_xcpt_ma_st;
	assign io_requestor_0_s2_xcpt_pf_ld = io_mem_s2_xcpt_pf_ld;
	assign io_requestor_0_s2_xcpt_pf_st = io_mem_s2_xcpt_pf_st;
	assign io_requestor_0_s2_xcpt_ae_ld = io_mem_s2_xcpt_ae_ld;
	assign io_requestor_0_s2_xcpt_ae_st = io_mem_s2_xcpt_ae_st;
	assign io_requestor_0_ordered = io_mem_ordered;
	assign io_requestor_0_perf_grant = io_mem_perf_grant;
	assign io_requestor_1_req_ready = io_requestor_0_req_ready & ~io_requestor_0_req_valid;
	assign io_requestor_1_s2_nack = io_mem_s2_nack & s2_id;
	assign io_requestor_1_resp_valid = io_mem_resp_valid & io_mem_resp_bits_tag[0];
	assign io_requestor_1_resp_bits_data_raw = io_mem_resp_bits_data_raw;
	assign io_mem_req_valid = io_requestor_0_req_valid | io_requestor_1_req_valid;
	assign io_mem_req_bits_addr = (io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr);
	assign io_mem_req_bits_tag = _GEN_1[6:0];
	assign io_mem_req_bits_cmd = (io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd);
	assign io_mem_req_bits_size = (io_requestor_0_req_valid ? io_requestor_0_req_bits_size : io_requestor_1_req_bits_size);
	assign io_mem_req_bits_signed = io_requestor_0_req_valid & io_requestor_0_req_bits_signed;
	assign io_mem_req_bits_dprv = (io_requestor_0_req_valid ? 2'h3 : 2'h0);
	assign io_mem_req_bits_no_xcpt = (io_requestor_0_req_valid ? 1'h0 : 1'h1);
	assign io_mem_s1_kill = (~s1_id ? io_requestor_0_s1_kill : io_requestor_1_s1_kill);
	assign io_mem_s1_data_data = (~s1_id ? io_requestor_0_s1_data_data : io_requestor_1_s1_data_data);
	assign io_mem_s1_data_mask = (~s1_id ? 4'h0 : io_requestor_1_s1_data_mask);
	always @(posedge clock) begin
		if (io_requestor_0_req_valid)
			s1_id <= 1'h0;
		else
			s1_id <= 1'h1;
		s2_id <= s1_id;
	end
endmodule
module OptimizationBarrier_21 (
	io_x,
	io_y
);
	input [2:0] io_x;
	output wire [2:0] io_y;
	assign io_y = io_x;
endmodule
module OptimizationBarrier_22 (
	io_x_ppn,
	io_x_d,
	io_x_a,
	io_x_u,
	io_x_x,
	io_x_w,
	io_x_r,
	io_y_ppn,
	io_y_d,
	io_y_a,
	io_y_u,
	io_y_x,
	io_y_w,
	io_y_r
);
	input [53:0] io_x_ppn;
	input io_x_d;
	input io_x_a;
	input io_x_u;
	input io_x_x;
	input io_x_w;
	input io_x_r;
	output wire [53:0] io_y_ppn;
	output wire io_y_d;
	output wire io_y_a;
	output wire io_y_u;
	output wire io_y_x;
	output wire io_y_w;
	output wire io_y_r;
	assign io_y_ppn = io_x_ppn;
	assign io_y_d = io_x_d;
	assign io_y_a = io_x_a;
	assign io_y_u = io_x_u;
	assign io_y_x = io_x_x;
	assign io_y_w = io_x_w;
	assign io_y_r = io_x_r;
endmodule
module PTW (
	clock,
	reset,
	io_requestor_0_status_debug,
	io_requestor_0_pmp_0_cfg_l,
	io_requestor_0_pmp_0_cfg_a,
	io_requestor_0_pmp_0_cfg_x,
	io_requestor_0_pmp_0_cfg_w,
	io_requestor_0_pmp_0_cfg_r,
	io_requestor_0_pmp_0_addr,
	io_requestor_0_pmp_0_mask,
	io_requestor_0_pmp_1_cfg_l,
	io_requestor_0_pmp_1_cfg_a,
	io_requestor_0_pmp_1_cfg_x,
	io_requestor_0_pmp_1_cfg_w,
	io_requestor_0_pmp_1_cfg_r,
	io_requestor_0_pmp_1_addr,
	io_requestor_0_pmp_1_mask,
	io_requestor_0_pmp_2_cfg_l,
	io_requestor_0_pmp_2_cfg_a,
	io_requestor_0_pmp_2_cfg_x,
	io_requestor_0_pmp_2_cfg_w,
	io_requestor_0_pmp_2_cfg_r,
	io_requestor_0_pmp_2_addr,
	io_requestor_0_pmp_2_mask,
	io_requestor_0_pmp_3_cfg_l,
	io_requestor_0_pmp_3_cfg_a,
	io_requestor_0_pmp_3_cfg_x,
	io_requestor_0_pmp_3_cfg_w,
	io_requestor_0_pmp_3_cfg_r,
	io_requestor_0_pmp_3_addr,
	io_requestor_0_pmp_3_mask,
	io_requestor_0_pmp_4_cfg_l,
	io_requestor_0_pmp_4_cfg_a,
	io_requestor_0_pmp_4_cfg_x,
	io_requestor_0_pmp_4_cfg_w,
	io_requestor_0_pmp_4_cfg_r,
	io_requestor_0_pmp_4_addr,
	io_requestor_0_pmp_4_mask,
	io_requestor_0_pmp_5_cfg_l,
	io_requestor_0_pmp_5_cfg_a,
	io_requestor_0_pmp_5_cfg_x,
	io_requestor_0_pmp_5_cfg_w,
	io_requestor_0_pmp_5_cfg_r,
	io_requestor_0_pmp_5_addr,
	io_requestor_0_pmp_5_mask,
	io_requestor_0_pmp_6_cfg_l,
	io_requestor_0_pmp_6_cfg_a,
	io_requestor_0_pmp_6_cfg_x,
	io_requestor_0_pmp_6_cfg_w,
	io_requestor_0_pmp_6_cfg_r,
	io_requestor_0_pmp_6_addr,
	io_requestor_0_pmp_6_mask,
	io_requestor_0_pmp_7_cfg_l,
	io_requestor_0_pmp_7_cfg_a,
	io_requestor_0_pmp_7_cfg_x,
	io_requestor_0_pmp_7_cfg_w,
	io_requestor_0_pmp_7_cfg_r,
	io_requestor_0_pmp_7_addr,
	io_requestor_0_pmp_7_mask,
	io_requestor_1_status_debug,
	io_requestor_1_pmp_0_cfg_l,
	io_requestor_1_pmp_0_cfg_a,
	io_requestor_1_pmp_0_cfg_x,
	io_requestor_1_pmp_0_cfg_w,
	io_requestor_1_pmp_0_cfg_r,
	io_requestor_1_pmp_0_addr,
	io_requestor_1_pmp_0_mask,
	io_requestor_1_pmp_1_cfg_l,
	io_requestor_1_pmp_1_cfg_a,
	io_requestor_1_pmp_1_cfg_x,
	io_requestor_1_pmp_1_cfg_w,
	io_requestor_1_pmp_1_cfg_r,
	io_requestor_1_pmp_1_addr,
	io_requestor_1_pmp_1_mask,
	io_requestor_1_pmp_2_cfg_l,
	io_requestor_1_pmp_2_cfg_a,
	io_requestor_1_pmp_2_cfg_x,
	io_requestor_1_pmp_2_cfg_w,
	io_requestor_1_pmp_2_cfg_r,
	io_requestor_1_pmp_2_addr,
	io_requestor_1_pmp_2_mask,
	io_requestor_1_pmp_3_cfg_l,
	io_requestor_1_pmp_3_cfg_a,
	io_requestor_1_pmp_3_cfg_x,
	io_requestor_1_pmp_3_cfg_w,
	io_requestor_1_pmp_3_cfg_r,
	io_requestor_1_pmp_3_addr,
	io_requestor_1_pmp_3_mask,
	io_requestor_1_pmp_4_cfg_l,
	io_requestor_1_pmp_4_cfg_a,
	io_requestor_1_pmp_4_cfg_x,
	io_requestor_1_pmp_4_cfg_w,
	io_requestor_1_pmp_4_cfg_r,
	io_requestor_1_pmp_4_addr,
	io_requestor_1_pmp_4_mask,
	io_requestor_1_pmp_5_cfg_l,
	io_requestor_1_pmp_5_cfg_a,
	io_requestor_1_pmp_5_cfg_x,
	io_requestor_1_pmp_5_cfg_w,
	io_requestor_1_pmp_5_cfg_r,
	io_requestor_1_pmp_5_addr,
	io_requestor_1_pmp_5_mask,
	io_requestor_1_pmp_6_cfg_l,
	io_requestor_1_pmp_6_cfg_a,
	io_requestor_1_pmp_6_cfg_x,
	io_requestor_1_pmp_6_cfg_w,
	io_requestor_1_pmp_6_cfg_r,
	io_requestor_1_pmp_6_addr,
	io_requestor_1_pmp_6_mask,
	io_requestor_1_pmp_7_cfg_l,
	io_requestor_1_pmp_7_cfg_a,
	io_requestor_1_pmp_7_cfg_x,
	io_requestor_1_pmp_7_cfg_w,
	io_requestor_1_pmp_7_cfg_r,
	io_requestor_1_pmp_7_addr,
	io_requestor_1_pmp_7_mask,
	io_requestor_1_customCSRs_csrs_0_value,
	io_dpath_status_debug,
	io_dpath_pmp_0_cfg_l,
	io_dpath_pmp_0_cfg_a,
	io_dpath_pmp_0_cfg_x,
	io_dpath_pmp_0_cfg_w,
	io_dpath_pmp_0_cfg_r,
	io_dpath_pmp_0_addr,
	io_dpath_pmp_0_mask,
	io_dpath_pmp_1_cfg_l,
	io_dpath_pmp_1_cfg_a,
	io_dpath_pmp_1_cfg_x,
	io_dpath_pmp_1_cfg_w,
	io_dpath_pmp_1_cfg_r,
	io_dpath_pmp_1_addr,
	io_dpath_pmp_1_mask,
	io_dpath_pmp_2_cfg_l,
	io_dpath_pmp_2_cfg_a,
	io_dpath_pmp_2_cfg_x,
	io_dpath_pmp_2_cfg_w,
	io_dpath_pmp_2_cfg_r,
	io_dpath_pmp_2_addr,
	io_dpath_pmp_2_mask,
	io_dpath_pmp_3_cfg_l,
	io_dpath_pmp_3_cfg_a,
	io_dpath_pmp_3_cfg_x,
	io_dpath_pmp_3_cfg_w,
	io_dpath_pmp_3_cfg_r,
	io_dpath_pmp_3_addr,
	io_dpath_pmp_3_mask,
	io_dpath_pmp_4_cfg_l,
	io_dpath_pmp_4_cfg_a,
	io_dpath_pmp_4_cfg_x,
	io_dpath_pmp_4_cfg_w,
	io_dpath_pmp_4_cfg_r,
	io_dpath_pmp_4_addr,
	io_dpath_pmp_4_mask,
	io_dpath_pmp_5_cfg_l,
	io_dpath_pmp_5_cfg_a,
	io_dpath_pmp_5_cfg_x,
	io_dpath_pmp_5_cfg_w,
	io_dpath_pmp_5_cfg_r,
	io_dpath_pmp_5_addr,
	io_dpath_pmp_5_mask,
	io_dpath_pmp_6_cfg_l,
	io_dpath_pmp_6_cfg_a,
	io_dpath_pmp_6_cfg_x,
	io_dpath_pmp_6_cfg_w,
	io_dpath_pmp_6_cfg_r,
	io_dpath_pmp_6_addr,
	io_dpath_pmp_6_mask,
	io_dpath_pmp_7_cfg_l,
	io_dpath_pmp_7_cfg_a,
	io_dpath_pmp_7_cfg_x,
	io_dpath_pmp_7_cfg_w,
	io_dpath_pmp_7_cfg_r,
	io_dpath_pmp_7_addr,
	io_dpath_pmp_7_mask,
	io_dpath_perf_l2hit,
	io_dpath_perf_pte_miss,
	io_dpath_perf_pte_hit,
	io_dpath_customCSRs_csrs_0_value
);
	input clock;
	input reset;
	output wire io_requestor_0_status_debug;
	output wire io_requestor_0_pmp_0_cfg_l;
	output wire [1:0] io_requestor_0_pmp_0_cfg_a;
	output wire io_requestor_0_pmp_0_cfg_x;
	output wire io_requestor_0_pmp_0_cfg_w;
	output wire io_requestor_0_pmp_0_cfg_r;
	output wire [29:0] io_requestor_0_pmp_0_addr;
	output wire [31:0] io_requestor_0_pmp_0_mask;
	output wire io_requestor_0_pmp_1_cfg_l;
	output wire [1:0] io_requestor_0_pmp_1_cfg_a;
	output wire io_requestor_0_pmp_1_cfg_x;
	output wire io_requestor_0_pmp_1_cfg_w;
	output wire io_requestor_0_pmp_1_cfg_r;
	output wire [29:0] io_requestor_0_pmp_1_addr;
	output wire [31:0] io_requestor_0_pmp_1_mask;
	output wire io_requestor_0_pmp_2_cfg_l;
	output wire [1:0] io_requestor_0_pmp_2_cfg_a;
	output wire io_requestor_0_pmp_2_cfg_x;
	output wire io_requestor_0_pmp_2_cfg_w;
	output wire io_requestor_0_pmp_2_cfg_r;
	output wire [29:0] io_requestor_0_pmp_2_addr;
	output wire [31:0] io_requestor_0_pmp_2_mask;
	output wire io_requestor_0_pmp_3_cfg_l;
	output wire [1:0] io_requestor_0_pmp_3_cfg_a;
	output wire io_requestor_0_pmp_3_cfg_x;
	output wire io_requestor_0_pmp_3_cfg_w;
	output wire io_requestor_0_pmp_3_cfg_r;
	output wire [29:0] io_requestor_0_pmp_3_addr;
	output wire [31:0] io_requestor_0_pmp_3_mask;
	output wire io_requestor_0_pmp_4_cfg_l;
	output wire [1:0] io_requestor_0_pmp_4_cfg_a;
	output wire io_requestor_0_pmp_4_cfg_x;
	output wire io_requestor_0_pmp_4_cfg_w;
	output wire io_requestor_0_pmp_4_cfg_r;
	output wire [29:0] io_requestor_0_pmp_4_addr;
	output wire [31:0] io_requestor_0_pmp_4_mask;
	output wire io_requestor_0_pmp_5_cfg_l;
	output wire [1:0] io_requestor_0_pmp_5_cfg_a;
	output wire io_requestor_0_pmp_5_cfg_x;
	output wire io_requestor_0_pmp_5_cfg_w;
	output wire io_requestor_0_pmp_5_cfg_r;
	output wire [29:0] io_requestor_0_pmp_5_addr;
	output wire [31:0] io_requestor_0_pmp_5_mask;
	output wire io_requestor_0_pmp_6_cfg_l;
	output wire [1:0] io_requestor_0_pmp_6_cfg_a;
	output wire io_requestor_0_pmp_6_cfg_x;
	output wire io_requestor_0_pmp_6_cfg_w;
	output wire io_requestor_0_pmp_6_cfg_r;
	output wire [29:0] io_requestor_0_pmp_6_addr;
	output wire [31:0] io_requestor_0_pmp_6_mask;
	output wire io_requestor_0_pmp_7_cfg_l;
	output wire [1:0] io_requestor_0_pmp_7_cfg_a;
	output wire io_requestor_0_pmp_7_cfg_x;
	output wire io_requestor_0_pmp_7_cfg_w;
	output wire io_requestor_0_pmp_7_cfg_r;
	output wire [29:0] io_requestor_0_pmp_7_addr;
	output wire [31:0] io_requestor_0_pmp_7_mask;
	output wire io_requestor_1_status_debug;
	output wire io_requestor_1_pmp_0_cfg_l;
	output wire [1:0] io_requestor_1_pmp_0_cfg_a;
	output wire io_requestor_1_pmp_0_cfg_x;
	output wire io_requestor_1_pmp_0_cfg_w;
	output wire io_requestor_1_pmp_0_cfg_r;
	output wire [29:0] io_requestor_1_pmp_0_addr;
	output wire [31:0] io_requestor_1_pmp_0_mask;
	output wire io_requestor_1_pmp_1_cfg_l;
	output wire [1:0] io_requestor_1_pmp_1_cfg_a;
	output wire io_requestor_1_pmp_1_cfg_x;
	output wire io_requestor_1_pmp_1_cfg_w;
	output wire io_requestor_1_pmp_1_cfg_r;
	output wire [29:0] io_requestor_1_pmp_1_addr;
	output wire [31:0] io_requestor_1_pmp_1_mask;
	output wire io_requestor_1_pmp_2_cfg_l;
	output wire [1:0] io_requestor_1_pmp_2_cfg_a;
	output wire io_requestor_1_pmp_2_cfg_x;
	output wire io_requestor_1_pmp_2_cfg_w;
	output wire io_requestor_1_pmp_2_cfg_r;
	output wire [29:0] io_requestor_1_pmp_2_addr;
	output wire [31:0] io_requestor_1_pmp_2_mask;
	output wire io_requestor_1_pmp_3_cfg_l;
	output wire [1:0] io_requestor_1_pmp_3_cfg_a;
	output wire io_requestor_1_pmp_3_cfg_x;
	output wire io_requestor_1_pmp_3_cfg_w;
	output wire io_requestor_1_pmp_3_cfg_r;
	output wire [29:0] io_requestor_1_pmp_3_addr;
	output wire [31:0] io_requestor_1_pmp_3_mask;
	output wire io_requestor_1_pmp_4_cfg_l;
	output wire [1:0] io_requestor_1_pmp_4_cfg_a;
	output wire io_requestor_1_pmp_4_cfg_x;
	output wire io_requestor_1_pmp_4_cfg_w;
	output wire io_requestor_1_pmp_4_cfg_r;
	output wire [29:0] io_requestor_1_pmp_4_addr;
	output wire [31:0] io_requestor_1_pmp_4_mask;
	output wire io_requestor_1_pmp_5_cfg_l;
	output wire [1:0] io_requestor_1_pmp_5_cfg_a;
	output wire io_requestor_1_pmp_5_cfg_x;
	output wire io_requestor_1_pmp_5_cfg_w;
	output wire io_requestor_1_pmp_5_cfg_r;
	output wire [29:0] io_requestor_1_pmp_5_addr;
	output wire [31:0] io_requestor_1_pmp_5_mask;
	output wire io_requestor_1_pmp_6_cfg_l;
	output wire [1:0] io_requestor_1_pmp_6_cfg_a;
	output wire io_requestor_1_pmp_6_cfg_x;
	output wire io_requestor_1_pmp_6_cfg_w;
	output wire io_requestor_1_pmp_6_cfg_r;
	output wire [29:0] io_requestor_1_pmp_6_addr;
	output wire [31:0] io_requestor_1_pmp_6_mask;
	output wire io_requestor_1_pmp_7_cfg_l;
	output wire [1:0] io_requestor_1_pmp_7_cfg_a;
	output wire io_requestor_1_pmp_7_cfg_x;
	output wire io_requestor_1_pmp_7_cfg_w;
	output wire io_requestor_1_pmp_7_cfg_r;
	output wire [29:0] io_requestor_1_pmp_7_addr;
	output wire [31:0] io_requestor_1_pmp_7_mask;
	output wire [31:0] io_requestor_1_customCSRs_csrs_0_value;
	input io_dpath_status_debug;
	input io_dpath_pmp_0_cfg_l;
	input [1:0] io_dpath_pmp_0_cfg_a;
	input io_dpath_pmp_0_cfg_x;
	input io_dpath_pmp_0_cfg_w;
	input io_dpath_pmp_0_cfg_r;
	input [29:0] io_dpath_pmp_0_addr;
	input [31:0] io_dpath_pmp_0_mask;
	input io_dpath_pmp_1_cfg_l;
	input [1:0] io_dpath_pmp_1_cfg_a;
	input io_dpath_pmp_1_cfg_x;
	input io_dpath_pmp_1_cfg_w;
	input io_dpath_pmp_1_cfg_r;
	input [29:0] io_dpath_pmp_1_addr;
	input [31:0] io_dpath_pmp_1_mask;
	input io_dpath_pmp_2_cfg_l;
	input [1:0] io_dpath_pmp_2_cfg_a;
	input io_dpath_pmp_2_cfg_x;
	input io_dpath_pmp_2_cfg_w;
	input io_dpath_pmp_2_cfg_r;
	input [29:0] io_dpath_pmp_2_addr;
	input [31:0] io_dpath_pmp_2_mask;
	input io_dpath_pmp_3_cfg_l;
	input [1:0] io_dpath_pmp_3_cfg_a;
	input io_dpath_pmp_3_cfg_x;
	input io_dpath_pmp_3_cfg_w;
	input io_dpath_pmp_3_cfg_r;
	input [29:0] io_dpath_pmp_3_addr;
	input [31:0] io_dpath_pmp_3_mask;
	input io_dpath_pmp_4_cfg_l;
	input [1:0] io_dpath_pmp_4_cfg_a;
	input io_dpath_pmp_4_cfg_x;
	input io_dpath_pmp_4_cfg_w;
	input io_dpath_pmp_4_cfg_r;
	input [29:0] io_dpath_pmp_4_addr;
	input [31:0] io_dpath_pmp_4_mask;
	input io_dpath_pmp_5_cfg_l;
	input [1:0] io_dpath_pmp_5_cfg_a;
	input io_dpath_pmp_5_cfg_x;
	input io_dpath_pmp_5_cfg_w;
	input io_dpath_pmp_5_cfg_r;
	input [29:0] io_dpath_pmp_5_addr;
	input [31:0] io_dpath_pmp_5_mask;
	input io_dpath_pmp_6_cfg_l;
	input [1:0] io_dpath_pmp_6_cfg_a;
	input io_dpath_pmp_6_cfg_x;
	input io_dpath_pmp_6_cfg_w;
	input io_dpath_pmp_6_cfg_r;
	input [29:0] io_dpath_pmp_6_addr;
	input [31:0] io_dpath_pmp_6_mask;
	input io_dpath_pmp_7_cfg_l;
	input [1:0] io_dpath_pmp_7_cfg_a;
	input io_dpath_pmp_7_cfg_x;
	input io_dpath_pmp_7_cfg_w;
	input io_dpath_pmp_7_cfg_r;
	input [29:0] io_dpath_pmp_7_addr;
	input [31:0] io_dpath_pmp_7_mask;
	output wire io_dpath_perf_l2hit;
	output wire io_dpath_perf_pte_miss;
	output wire io_dpath_perf_pte_hit;
	input [31:0] io_dpath_customCSRs_csrs_0_value;
	wire l2_tlb_ram_RW0_clk;
	wire [36:0] l2_tlb_ram_RW0_wdata_0;
	wire [2:0] state_barrier_io_x;
	wire [2:0] state_barrier_io_y;
	wire [53:0] r_pte_barrier_io_x_ppn;
	wire r_pte_barrier_io_x_d;
	wire r_pte_barrier_io_x_a;
	wire r_pte_barrier_io_x_u;
	wire r_pte_barrier_io_x_x;
	wire r_pte_barrier_io_x_w;
	wire r_pte_barrier_io_x_r;
	wire [53:0] r_pte_barrier_io_y_ppn;
	wire r_pte_barrier_io_y_d;
	wire r_pte_barrier_io_y_a;
	wire r_pte_barrier_io_y_u;
	wire r_pte_barrier_io_y_x;
	wire r_pte_barrier_io_y_w;
	wire r_pte_barrier_io_y_r;
	reg [2:0] state;
	reg [53:0] r_pte_ppn;
	reg r_pte_d;
	reg r_pte_a;
	reg r_pte_u;
	reg r_pte_x;
	reg r_pte_w;
	reg r_pte_r;
	wire [19:0] entry_ppn = r_pte_ppn[19:0];
	wire [35:0] _T_132 = {10'h000, entry_ppn, r_pte_d, r_pte_a, r_pte_u, r_pte_x, r_pte_w, r_pte_r};
	wire _T_133 = ^_T_132;
	wire [65:0] _pmaPgLevelHomogeneous_T = {r_pte_ppn, 12'h000};
	wire [65:0] _pmaPgLevelHomogeneous_T_1 = _pmaPgLevelHomogeneous_T ^ 66'h0000000000c000000;
	wire [66:0] _pmaPgLevelHomogeneous_T_2 = {1'b0, $signed(_pmaPgLevelHomogeneous_T_1)};
	wire [66:0] _pmaPgLevelHomogeneous_T_4 = $signed(_pmaPgLevelHomogeneous_T_2) & -67'sh00000000004000000;
	wire pmaPgLevelHomogeneous_0 = $signed(_pmaPgLevelHomogeneous_T_4) == 67'sh00000000000000000;
	wire [66:0] _pmaPgLevelHomogeneous_T_12 = {1'b0, $signed(_pmaPgLevelHomogeneous_T)};
	wire [66:0] _pmaPgLevelHomogeneous_T_14 = $signed(_pmaPgLevelHomogeneous_T_12) & -67'sh00000000000005000;
	wire _pmaPgLevelHomogeneous_T_15 = $signed(_pmaPgLevelHomogeneous_T_14) == 67'sh00000000000000000;
	wire [65:0] _pmaPgLevelHomogeneous_T_16 = _pmaPgLevelHomogeneous_T ^ 66'h00000000000003000;
	wire [66:0] _pmaPgLevelHomogeneous_T_17 = {1'b0, $signed(_pmaPgLevelHomogeneous_T_16)};
	wire [66:0] _pmaPgLevelHomogeneous_T_19 = $signed(_pmaPgLevelHomogeneous_T_17) & -67'sh00000000000001000;
	wire _pmaPgLevelHomogeneous_T_20 = $signed(_pmaPgLevelHomogeneous_T_19) == 67'sh00000000000000000;
	wire [65:0] _pmaPgLevelHomogeneous_T_21 = _pmaPgLevelHomogeneous_T ^ 66'h00000000000010000;
	wire [66:0] _pmaPgLevelHomogeneous_T_22 = {1'b0, $signed(_pmaPgLevelHomogeneous_T_21)};
	wire [66:0] _pmaPgLevelHomogeneous_T_24 = $signed(_pmaPgLevelHomogeneous_T_22) & -67'sh00000000000010000;
	wire _pmaPgLevelHomogeneous_T_25 = $signed(_pmaPgLevelHomogeneous_T_24) == 67'sh00000000000000000;
	wire [65:0] _pmaPgLevelHomogeneous_T_26 = _pmaPgLevelHomogeneous_T ^ 66'h00000000000020000;
	wire [66:0] _pmaPgLevelHomogeneous_T_27 = {1'b0, $signed(_pmaPgLevelHomogeneous_T_26)};
	wire [66:0] _pmaPgLevelHomogeneous_T_29 = $signed(_pmaPgLevelHomogeneous_T_27) & -67'sh00000000000010000;
	wire _pmaPgLevelHomogeneous_T_30 = $signed(_pmaPgLevelHomogeneous_T_29) == 67'sh00000000000000000;
	wire [65:0] _pmaPgLevelHomogeneous_T_31 = _pmaPgLevelHomogeneous_T ^ 66'h00000000000100000;
	wire [66:0] _pmaPgLevelHomogeneous_T_32 = {1'b0, $signed(_pmaPgLevelHomogeneous_T_31)};
	wire [66:0] _pmaPgLevelHomogeneous_T_34 = $signed(_pmaPgLevelHomogeneous_T_32) & -67'sh00000000000011000;
	wire _pmaPgLevelHomogeneous_T_35 = $signed(_pmaPgLevelHomogeneous_T_34) == 67'sh00000000000000000;
	wire [65:0] _pmaPgLevelHomogeneous_T_36 = _pmaPgLevelHomogeneous_T ^ 66'h00000000002000000;
	wire [66:0] _pmaPgLevelHomogeneous_T_37 = {1'b0, $signed(_pmaPgLevelHomogeneous_T_36)};
	wire [66:0] _pmaPgLevelHomogeneous_T_39 = $signed(_pmaPgLevelHomogeneous_T_37) & -67'sh00000000000010000;
	wire _pmaPgLevelHomogeneous_T_40 = $signed(_pmaPgLevelHomogeneous_T_39) == 67'sh00000000000000000;
	wire [65:0] _pmaPgLevelHomogeneous_T_46 = _pmaPgLevelHomogeneous_T ^ 66'h00000000010000000;
	wire [66:0] _pmaPgLevelHomogeneous_T_47 = {1'b0, $signed(_pmaPgLevelHomogeneous_T_46)};
	wire [66:0] _pmaPgLevelHomogeneous_T_49 = $signed(_pmaPgLevelHomogeneous_T_47) & -67'sh00000000000001000;
	wire _pmaPgLevelHomogeneous_T_50 = $signed(_pmaPgLevelHomogeneous_T_49) == 67'sh00000000000000000;
	wire [65:0] _pmaPgLevelHomogeneous_T_51 = _pmaPgLevelHomogeneous_T ^ 66'h00000000054000000;
	wire [66:0] _pmaPgLevelHomogeneous_T_52 = {1'b0, $signed(_pmaPgLevelHomogeneous_T_51)};
	wire [66:0] _pmaPgLevelHomogeneous_T_54 = $signed(_pmaPgLevelHomogeneous_T_52) & -67'sh00000000000001000;
	wire _pmaPgLevelHomogeneous_T_55 = $signed(_pmaPgLevelHomogeneous_T_54) == 67'sh00000000000000000;
	wire [65:0] _pmaPgLevelHomogeneous_T_56 = _pmaPgLevelHomogeneous_T ^ 66'h00000000080000000;
	wire [66:0] _pmaPgLevelHomogeneous_T_57 = {1'b0, $signed(_pmaPgLevelHomogeneous_T_56)};
	wire [66:0] _pmaPgLevelHomogeneous_T_59 = $signed(_pmaPgLevelHomogeneous_T_57) & -67'sh00000000000004000;
	wire _pmaPgLevelHomogeneous_T_60 = $signed(_pmaPgLevelHomogeneous_T_59) == 67'sh00000000000000000;
	wire pmaPgLevelHomogeneous_1 = ((((((((_pmaPgLevelHomogeneous_T_15 | _pmaPgLevelHomogeneous_T_20) | _pmaPgLevelHomogeneous_T_25) | _pmaPgLevelHomogeneous_T_30) | _pmaPgLevelHomogeneous_T_35) | _pmaPgLevelHomogeneous_T_40) | pmaPgLevelHomogeneous_0) | _pmaPgLevelHomogeneous_T_50) | _pmaPgLevelHomogeneous_T_55) | _pmaPgLevelHomogeneous_T_60;
	wire pmpHomogeneous_maskHomogeneous = io_dpath_pmp_0_mask[11];
	wire [31:0] _pmpHomogeneous_T_2 = {io_dpath_pmp_0_addr, 2'h0};
	wire [31:0] _pmpHomogeneous_T_3 = ~_pmpHomogeneous_T_2;
	wire [31:0] _pmpHomogeneous_T_4 = _pmpHomogeneous_T_3 | 32'h00000003;
	wire [31:0] _pmpHomogeneous_T_5 = ~_pmpHomogeneous_T_4;
	wire [65:0] _GEN_94 = {34'd0, _pmpHomogeneous_T_5};
	wire [65:0] _pmpHomogeneous_T_6 = _pmaPgLevelHomogeneous_T ^ _GEN_94;
	wire _pmpHomogeneous_T_18 = pmpHomogeneous_maskHomogeneous | (_pmpHomogeneous_T_6[65:12] != 54'h00000000000000);
	wire pmpHomogeneous_beginsAfterUpper = ~(_pmaPgLevelHomogeneous_T < _GEN_94);
	wire [65:0] _pmpHomogeneous_endsBeforeLower_T = _pmaPgLevelHomogeneous_T & 66'h000000000fffff000;
	wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_5 = _pmpHomogeneous_T_5 & 32'hfffff000;
	wire [65:0] _GEN_97 = {34'd0, _pmpHomogeneous_endsBeforeUpper_T_5};
	wire pmpHomogeneous_endsBeforeUpper = _pmpHomogeneous_endsBeforeLower_T < _GEN_97;
	wire _pmpHomogeneous_T_23 = pmpHomogeneous_beginsAfterUpper | pmpHomogeneous_endsBeforeUpper;
	wire _pmpHomogeneous_T_25 = (io_dpath_pmp_0_cfg_a[1] ? _pmpHomogeneous_T_18 : ~io_dpath_pmp_0_cfg_a[0] | _pmpHomogeneous_T_23);
	wire pmpHomogeneous_maskHomogeneous_1 = io_dpath_pmp_1_mask[11];
	wire [31:0] _pmpHomogeneous_T_28 = {io_dpath_pmp_1_addr, 2'h0};
	wire [31:0] _pmpHomogeneous_T_29 = ~_pmpHomogeneous_T_28;
	wire [31:0] _pmpHomogeneous_T_30 = _pmpHomogeneous_T_29 | 32'h00000003;
	wire [31:0] _pmpHomogeneous_T_31 = ~_pmpHomogeneous_T_30;
	wire [65:0] _GEN_98 = {34'd0, _pmpHomogeneous_T_31};
	wire [65:0] _pmpHomogeneous_T_32 = _pmaPgLevelHomogeneous_T ^ _GEN_98;
	wire _pmpHomogeneous_T_44 = pmpHomogeneous_maskHomogeneous_1 | (_pmpHomogeneous_T_32[65:12] != 54'h00000000000000);
	wire pmpHomogeneous_beginsAfterUpper_1 = ~(_pmaPgLevelHomogeneous_T < _GEN_98);
	wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_11 = _pmpHomogeneous_T_31 & 32'hfffff000;
	wire [65:0] _GEN_103 = {34'd0, _pmpHomogeneous_endsBeforeUpper_T_11};
	wire pmpHomogeneous_endsBeforeUpper_1 = _pmpHomogeneous_endsBeforeLower_T < _GEN_103;
	wire _pmpHomogeneous_T_49 = (pmpHomogeneous_endsBeforeUpper | pmpHomogeneous_beginsAfterUpper_1) | (pmpHomogeneous_beginsAfterUpper & pmpHomogeneous_endsBeforeUpper_1);
	wire _pmpHomogeneous_T_51 = (io_dpath_pmp_1_cfg_a[1] ? _pmpHomogeneous_T_44 : ~io_dpath_pmp_1_cfg_a[0] | _pmpHomogeneous_T_49);
	wire pmpHomogeneous_maskHomogeneous_2 = io_dpath_pmp_2_mask[11];
	wire [31:0] _pmpHomogeneous_T_54 = {io_dpath_pmp_2_addr, 2'h0};
	wire [31:0] _pmpHomogeneous_T_55 = ~_pmpHomogeneous_T_54;
	wire [31:0] _pmpHomogeneous_T_56 = _pmpHomogeneous_T_55 | 32'h00000003;
	wire [31:0] _pmpHomogeneous_T_57 = ~_pmpHomogeneous_T_56;
	wire [65:0] _GEN_104 = {34'd0, _pmpHomogeneous_T_57};
	wire [65:0] _pmpHomogeneous_T_58 = _pmaPgLevelHomogeneous_T ^ _GEN_104;
	wire _pmpHomogeneous_T_70 = pmpHomogeneous_maskHomogeneous_2 | (_pmpHomogeneous_T_58[65:12] != 54'h00000000000000);
	wire pmpHomogeneous_beginsAfterUpper_2 = ~(_pmaPgLevelHomogeneous_T < _GEN_104);
	wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_17 = _pmpHomogeneous_T_57 & 32'hfffff000;
	wire [65:0] _GEN_109 = {34'd0, _pmpHomogeneous_endsBeforeUpper_T_17};
	wire pmpHomogeneous_endsBeforeUpper_2 = _pmpHomogeneous_endsBeforeLower_T < _GEN_109;
	wire _pmpHomogeneous_T_75 = (pmpHomogeneous_endsBeforeUpper_1 | pmpHomogeneous_beginsAfterUpper_2) | (pmpHomogeneous_beginsAfterUpper_1 & pmpHomogeneous_endsBeforeUpper_2);
	wire _pmpHomogeneous_T_77 = (io_dpath_pmp_2_cfg_a[1] ? _pmpHomogeneous_T_70 : ~io_dpath_pmp_2_cfg_a[0] | _pmpHomogeneous_T_75);
	wire pmpHomogeneous_maskHomogeneous_3 = io_dpath_pmp_3_mask[11];
	wire [31:0] _pmpHomogeneous_T_80 = {io_dpath_pmp_3_addr, 2'h0};
	wire [31:0] _pmpHomogeneous_T_81 = ~_pmpHomogeneous_T_80;
	wire [31:0] _pmpHomogeneous_T_82 = _pmpHomogeneous_T_81 | 32'h00000003;
	wire [31:0] _pmpHomogeneous_T_83 = ~_pmpHomogeneous_T_82;
	wire [65:0] _GEN_110 = {34'd0, _pmpHomogeneous_T_83};
	wire [65:0] _pmpHomogeneous_T_84 = _pmaPgLevelHomogeneous_T ^ _GEN_110;
	wire _pmpHomogeneous_T_96 = pmpHomogeneous_maskHomogeneous_3 | (_pmpHomogeneous_T_84[65:12] != 54'h00000000000000);
	wire pmpHomogeneous_beginsAfterUpper_3 = ~(_pmaPgLevelHomogeneous_T < _GEN_110);
	wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_23 = _pmpHomogeneous_T_83 & 32'hfffff000;
	wire [65:0] _GEN_115 = {34'd0, _pmpHomogeneous_endsBeforeUpper_T_23};
	wire pmpHomogeneous_endsBeforeUpper_3 = _pmpHomogeneous_endsBeforeLower_T < _GEN_115;
	wire _pmpHomogeneous_T_101 = (pmpHomogeneous_endsBeforeUpper_2 | pmpHomogeneous_beginsAfterUpper_3) | (pmpHomogeneous_beginsAfterUpper_2 & pmpHomogeneous_endsBeforeUpper_3);
	wire _pmpHomogeneous_T_103 = (io_dpath_pmp_3_cfg_a[1] ? _pmpHomogeneous_T_96 : ~io_dpath_pmp_3_cfg_a[0] | _pmpHomogeneous_T_101);
	wire pmpHomogeneous_maskHomogeneous_4 = io_dpath_pmp_4_mask[11];
	wire [31:0] _pmpHomogeneous_T_106 = {io_dpath_pmp_4_addr, 2'h0};
	wire [31:0] _pmpHomogeneous_T_107 = ~_pmpHomogeneous_T_106;
	wire [31:0] _pmpHomogeneous_T_108 = _pmpHomogeneous_T_107 | 32'h00000003;
	wire [31:0] _pmpHomogeneous_T_109 = ~_pmpHomogeneous_T_108;
	wire [65:0] _GEN_116 = {34'd0, _pmpHomogeneous_T_109};
	wire [65:0] _pmpHomogeneous_T_110 = _pmaPgLevelHomogeneous_T ^ _GEN_116;
	wire _pmpHomogeneous_T_122 = pmpHomogeneous_maskHomogeneous_4 | (_pmpHomogeneous_T_110[65:12] != 54'h00000000000000);
	wire pmpHomogeneous_beginsAfterUpper_4 = ~(_pmaPgLevelHomogeneous_T < _GEN_116);
	wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_29 = _pmpHomogeneous_T_109 & 32'hfffff000;
	wire [65:0] _GEN_121 = {34'd0, _pmpHomogeneous_endsBeforeUpper_T_29};
	wire pmpHomogeneous_endsBeforeUpper_4 = _pmpHomogeneous_endsBeforeLower_T < _GEN_121;
	wire _pmpHomogeneous_T_127 = (pmpHomogeneous_endsBeforeUpper_3 | pmpHomogeneous_beginsAfterUpper_4) | (pmpHomogeneous_beginsAfterUpper_3 & pmpHomogeneous_endsBeforeUpper_4);
	wire _pmpHomogeneous_T_129 = (io_dpath_pmp_4_cfg_a[1] ? _pmpHomogeneous_T_122 : ~io_dpath_pmp_4_cfg_a[0] | _pmpHomogeneous_T_127);
	wire pmpHomogeneous_maskHomogeneous_5 = io_dpath_pmp_5_mask[11];
	wire [31:0] _pmpHomogeneous_T_132 = {io_dpath_pmp_5_addr, 2'h0};
	wire [31:0] _pmpHomogeneous_T_133 = ~_pmpHomogeneous_T_132;
	wire [31:0] _pmpHomogeneous_T_134 = _pmpHomogeneous_T_133 | 32'h00000003;
	wire [31:0] _pmpHomogeneous_T_135 = ~_pmpHomogeneous_T_134;
	wire [65:0] _GEN_122 = {34'd0, _pmpHomogeneous_T_135};
	wire [65:0] _pmpHomogeneous_T_136 = _pmaPgLevelHomogeneous_T ^ _GEN_122;
	wire _pmpHomogeneous_T_148 = pmpHomogeneous_maskHomogeneous_5 | (_pmpHomogeneous_T_136[65:12] != 54'h00000000000000);
	wire pmpHomogeneous_beginsAfterUpper_5 = ~(_pmaPgLevelHomogeneous_T < _GEN_122);
	wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_35 = _pmpHomogeneous_T_135 & 32'hfffff000;
	wire [65:0] _GEN_127 = {34'd0, _pmpHomogeneous_endsBeforeUpper_T_35};
	wire pmpHomogeneous_endsBeforeUpper_5 = _pmpHomogeneous_endsBeforeLower_T < _GEN_127;
	wire _pmpHomogeneous_T_153 = (pmpHomogeneous_endsBeforeUpper_4 | pmpHomogeneous_beginsAfterUpper_5) | (pmpHomogeneous_beginsAfterUpper_4 & pmpHomogeneous_endsBeforeUpper_5);
	wire _pmpHomogeneous_T_155 = (io_dpath_pmp_5_cfg_a[1] ? _pmpHomogeneous_T_148 : ~io_dpath_pmp_5_cfg_a[0] | _pmpHomogeneous_T_153);
	wire pmpHomogeneous_maskHomogeneous_6 = io_dpath_pmp_6_mask[11];
	wire [31:0] _pmpHomogeneous_T_158 = {io_dpath_pmp_6_addr, 2'h0};
	wire [31:0] _pmpHomogeneous_T_159 = ~_pmpHomogeneous_T_158;
	wire [31:0] _pmpHomogeneous_T_160 = _pmpHomogeneous_T_159 | 32'h00000003;
	wire [31:0] _pmpHomogeneous_T_161 = ~_pmpHomogeneous_T_160;
	wire [65:0] _GEN_128 = {34'd0, _pmpHomogeneous_T_161};
	wire [65:0] _pmpHomogeneous_T_162 = _pmaPgLevelHomogeneous_T ^ _GEN_128;
	wire _pmpHomogeneous_T_174 = pmpHomogeneous_maskHomogeneous_6 | (_pmpHomogeneous_T_162[65:12] != 54'h00000000000000);
	wire pmpHomogeneous_beginsAfterUpper_6 = ~(_pmaPgLevelHomogeneous_T < _GEN_128);
	wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_41 = _pmpHomogeneous_T_161 & 32'hfffff000;
	wire [65:0] _GEN_133 = {34'd0, _pmpHomogeneous_endsBeforeUpper_T_41};
	wire pmpHomogeneous_endsBeforeUpper_6 = _pmpHomogeneous_endsBeforeLower_T < _GEN_133;
	wire _pmpHomogeneous_T_179 = (pmpHomogeneous_endsBeforeUpper_5 | pmpHomogeneous_beginsAfterUpper_6) | (pmpHomogeneous_beginsAfterUpper_5 & pmpHomogeneous_endsBeforeUpper_6);
	wire _pmpHomogeneous_T_181 = (io_dpath_pmp_6_cfg_a[1] ? _pmpHomogeneous_T_174 : ~io_dpath_pmp_6_cfg_a[0] | _pmpHomogeneous_T_179);
	wire pmpHomogeneous_maskHomogeneous_7 = io_dpath_pmp_7_mask[11];
	wire [31:0] _pmpHomogeneous_T_184 = {io_dpath_pmp_7_addr, 2'h0};
	wire [31:0] _pmpHomogeneous_T_185 = ~_pmpHomogeneous_T_184;
	wire [31:0] _pmpHomogeneous_T_186 = _pmpHomogeneous_T_185 | 32'h00000003;
	wire [31:0] _pmpHomogeneous_T_187 = ~_pmpHomogeneous_T_186;
	wire [65:0] _GEN_134 = {34'd0, _pmpHomogeneous_T_187};
	wire [65:0] _pmpHomogeneous_T_188 = _pmaPgLevelHomogeneous_T ^ _GEN_134;
	wire _pmpHomogeneous_T_200 = pmpHomogeneous_maskHomogeneous_7 | (_pmpHomogeneous_T_188[65:12] != 54'h00000000000000);
	wire pmpHomogeneous_beginsAfterUpper_7 = ~(_pmaPgLevelHomogeneous_T < _GEN_134);
	wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_47 = _pmpHomogeneous_T_187 & 32'hfffff000;
	wire [65:0] _GEN_139 = {34'd0, _pmpHomogeneous_endsBeforeUpper_T_47};
	wire pmpHomogeneous_endsBeforeUpper_7 = _pmpHomogeneous_endsBeforeLower_T < _GEN_139;
	wire _pmpHomogeneous_T_205 = (pmpHomogeneous_endsBeforeUpper_6 | pmpHomogeneous_beginsAfterUpper_7) | (pmpHomogeneous_beginsAfterUpper_6 & pmpHomogeneous_endsBeforeUpper_7);
	wire _pmpHomogeneous_T_207 = (io_dpath_pmp_7_cfg_a[1] ? _pmpHomogeneous_T_200 : ~io_dpath_pmp_7_cfg_a[0] | _pmpHomogeneous_T_205);
	wire pmpHomogeneous = ((((((_pmpHomogeneous_T_25 & _pmpHomogeneous_T_51) & _pmpHomogeneous_T_77) & _pmpHomogeneous_T_103) & _pmpHomogeneous_T_129) & _pmpHomogeneous_T_155) & _pmpHomogeneous_T_181) & _pmpHomogeneous_T_207;
	wire homogeneous = pmaPgLevelHomogeneous_1 & pmpHomogeneous;
	wire _T_199 = ~homogeneous;
	wire [2:0] _GEN_2183 = (3'h7 == state ? 3'h0 : state);
	wire [2:0] _GEN_2188 = (3'h4 == state ? 3'h5 : _GEN_2183);
	wire [2:0] _GEN_2195 = (3'h2 == state ? 3'h4 : _GEN_2188);
	wire [2:0] _GEN_2207 = (3'h1 == state ? 3'h1 : _GEN_2195);
	wire [53:0] pte_2_ppn = {r_pte_ppn[53:10], 10'h000};
	l2_tlb_ram l2_tlb_ram(
		.RW0_clk(l2_tlb_ram_RW0_clk),
		.RW0_wdata_0(l2_tlb_ram_RW0_wdata_0)
	);
	OptimizationBarrier_21 state_barrier(
		.io_x(state_barrier_io_x),
		.io_y(state_barrier_io_y)
	);
	OptimizationBarrier_22 r_pte_barrier(
		.io_x_ppn(r_pte_barrier_io_x_ppn),
		.io_x_d(r_pte_barrier_io_x_d),
		.io_x_a(r_pte_barrier_io_x_a),
		.io_x_u(r_pte_barrier_io_x_u),
		.io_x_x(r_pte_barrier_io_x_x),
		.io_x_w(r_pte_barrier_io_x_w),
		.io_x_r(r_pte_barrier_io_x_r),
		.io_y_ppn(r_pte_barrier_io_y_ppn),
		.io_y_d(r_pte_barrier_io_y_d),
		.io_y_a(r_pte_barrier_io_y_a),
		.io_y_u(r_pte_barrier_io_y_u),
		.io_y_x(r_pte_barrier_io_y_x),
		.io_y_w(r_pte_barrier_io_y_w),
		.io_y_r(r_pte_barrier_io_y_r)
	);
	assign io_requestor_0_status_debug = io_dpath_status_debug;
	assign io_requestor_0_pmp_0_cfg_l = io_dpath_pmp_0_cfg_l;
	assign io_requestor_0_pmp_0_cfg_a = io_dpath_pmp_0_cfg_a;
	assign io_requestor_0_pmp_0_cfg_x = io_dpath_pmp_0_cfg_x;
	assign io_requestor_0_pmp_0_cfg_w = io_dpath_pmp_0_cfg_w;
	assign io_requestor_0_pmp_0_cfg_r = io_dpath_pmp_0_cfg_r;
	assign io_requestor_0_pmp_0_addr = io_dpath_pmp_0_addr;
	assign io_requestor_0_pmp_0_mask = io_dpath_pmp_0_mask;
	assign io_requestor_0_pmp_1_cfg_l = io_dpath_pmp_1_cfg_l;
	assign io_requestor_0_pmp_1_cfg_a = io_dpath_pmp_1_cfg_a;
	assign io_requestor_0_pmp_1_cfg_x = io_dpath_pmp_1_cfg_x;
	assign io_requestor_0_pmp_1_cfg_w = io_dpath_pmp_1_cfg_w;
	assign io_requestor_0_pmp_1_cfg_r = io_dpath_pmp_1_cfg_r;
	assign io_requestor_0_pmp_1_addr = io_dpath_pmp_1_addr;
	assign io_requestor_0_pmp_1_mask = io_dpath_pmp_1_mask;
	assign io_requestor_0_pmp_2_cfg_l = io_dpath_pmp_2_cfg_l;
	assign io_requestor_0_pmp_2_cfg_a = io_dpath_pmp_2_cfg_a;
	assign io_requestor_0_pmp_2_cfg_x = io_dpath_pmp_2_cfg_x;
	assign io_requestor_0_pmp_2_cfg_w = io_dpath_pmp_2_cfg_w;
	assign io_requestor_0_pmp_2_cfg_r = io_dpath_pmp_2_cfg_r;
	assign io_requestor_0_pmp_2_addr = io_dpath_pmp_2_addr;
	assign io_requestor_0_pmp_2_mask = io_dpath_pmp_2_mask;
	assign io_requestor_0_pmp_3_cfg_l = io_dpath_pmp_3_cfg_l;
	assign io_requestor_0_pmp_3_cfg_a = io_dpath_pmp_3_cfg_a;
	assign io_requestor_0_pmp_3_cfg_x = io_dpath_pmp_3_cfg_x;
	assign io_requestor_0_pmp_3_cfg_w = io_dpath_pmp_3_cfg_w;
	assign io_requestor_0_pmp_3_cfg_r = io_dpath_pmp_3_cfg_r;
	assign io_requestor_0_pmp_3_addr = io_dpath_pmp_3_addr;
	assign io_requestor_0_pmp_3_mask = io_dpath_pmp_3_mask;
	assign io_requestor_0_pmp_4_cfg_l = io_dpath_pmp_4_cfg_l;
	assign io_requestor_0_pmp_4_cfg_a = io_dpath_pmp_4_cfg_a;
	assign io_requestor_0_pmp_4_cfg_x = io_dpath_pmp_4_cfg_x;
	assign io_requestor_0_pmp_4_cfg_w = io_dpath_pmp_4_cfg_w;
	assign io_requestor_0_pmp_4_cfg_r = io_dpath_pmp_4_cfg_r;
	assign io_requestor_0_pmp_4_addr = io_dpath_pmp_4_addr;
	assign io_requestor_0_pmp_4_mask = io_dpath_pmp_4_mask;
	assign io_requestor_0_pmp_5_cfg_l = io_dpath_pmp_5_cfg_l;
	assign io_requestor_0_pmp_5_cfg_a = io_dpath_pmp_5_cfg_a;
	assign io_requestor_0_pmp_5_cfg_x = io_dpath_pmp_5_cfg_x;
	assign io_requestor_0_pmp_5_cfg_w = io_dpath_pmp_5_cfg_w;
	assign io_requestor_0_pmp_5_cfg_r = io_dpath_pmp_5_cfg_r;
	assign io_requestor_0_pmp_5_addr = io_dpath_pmp_5_addr;
	assign io_requestor_0_pmp_5_mask = io_dpath_pmp_5_mask;
	assign io_requestor_0_pmp_6_cfg_l = io_dpath_pmp_6_cfg_l;
	assign io_requestor_0_pmp_6_cfg_a = io_dpath_pmp_6_cfg_a;
	assign io_requestor_0_pmp_6_cfg_x = io_dpath_pmp_6_cfg_x;
	assign io_requestor_0_pmp_6_cfg_w = io_dpath_pmp_6_cfg_w;
	assign io_requestor_0_pmp_6_cfg_r = io_dpath_pmp_6_cfg_r;
	assign io_requestor_0_pmp_6_addr = io_dpath_pmp_6_addr;
	assign io_requestor_0_pmp_6_mask = io_dpath_pmp_6_mask;
	assign io_requestor_0_pmp_7_cfg_l = io_dpath_pmp_7_cfg_l;
	assign io_requestor_0_pmp_7_cfg_a = io_dpath_pmp_7_cfg_a;
	assign io_requestor_0_pmp_7_cfg_x = io_dpath_pmp_7_cfg_x;
	assign io_requestor_0_pmp_7_cfg_w = io_dpath_pmp_7_cfg_w;
	assign io_requestor_0_pmp_7_cfg_r = io_dpath_pmp_7_cfg_r;
	assign io_requestor_0_pmp_7_addr = io_dpath_pmp_7_addr;
	assign io_requestor_0_pmp_7_mask = io_dpath_pmp_7_mask;
	assign io_requestor_1_status_debug = io_dpath_status_debug;
	assign io_requestor_1_pmp_0_cfg_l = io_dpath_pmp_0_cfg_l;
	assign io_requestor_1_pmp_0_cfg_a = io_dpath_pmp_0_cfg_a;
	assign io_requestor_1_pmp_0_cfg_x = io_dpath_pmp_0_cfg_x;
	assign io_requestor_1_pmp_0_cfg_w = io_dpath_pmp_0_cfg_w;
	assign io_requestor_1_pmp_0_cfg_r = io_dpath_pmp_0_cfg_r;
	assign io_requestor_1_pmp_0_addr = io_dpath_pmp_0_addr;
	assign io_requestor_1_pmp_0_mask = io_dpath_pmp_0_mask;
	assign io_requestor_1_pmp_1_cfg_l = io_dpath_pmp_1_cfg_l;
	assign io_requestor_1_pmp_1_cfg_a = io_dpath_pmp_1_cfg_a;
	assign io_requestor_1_pmp_1_cfg_x = io_dpath_pmp_1_cfg_x;
	assign io_requestor_1_pmp_1_cfg_w = io_dpath_pmp_1_cfg_w;
	assign io_requestor_1_pmp_1_cfg_r = io_dpath_pmp_1_cfg_r;
	assign io_requestor_1_pmp_1_addr = io_dpath_pmp_1_addr;
	assign io_requestor_1_pmp_1_mask = io_dpath_pmp_1_mask;
	assign io_requestor_1_pmp_2_cfg_l = io_dpath_pmp_2_cfg_l;
	assign io_requestor_1_pmp_2_cfg_a = io_dpath_pmp_2_cfg_a;
	assign io_requestor_1_pmp_2_cfg_x = io_dpath_pmp_2_cfg_x;
	assign io_requestor_1_pmp_2_cfg_w = io_dpath_pmp_2_cfg_w;
	assign io_requestor_1_pmp_2_cfg_r = io_dpath_pmp_2_cfg_r;
	assign io_requestor_1_pmp_2_addr = io_dpath_pmp_2_addr;
	assign io_requestor_1_pmp_2_mask = io_dpath_pmp_2_mask;
	assign io_requestor_1_pmp_3_cfg_l = io_dpath_pmp_3_cfg_l;
	assign io_requestor_1_pmp_3_cfg_a = io_dpath_pmp_3_cfg_a;
	assign io_requestor_1_pmp_3_cfg_x = io_dpath_pmp_3_cfg_x;
	assign io_requestor_1_pmp_3_cfg_w = io_dpath_pmp_3_cfg_w;
	assign io_requestor_1_pmp_3_cfg_r = io_dpath_pmp_3_cfg_r;
	assign io_requestor_1_pmp_3_addr = io_dpath_pmp_3_addr;
	assign io_requestor_1_pmp_3_mask = io_dpath_pmp_3_mask;
	assign io_requestor_1_pmp_4_cfg_l = io_dpath_pmp_4_cfg_l;
	assign io_requestor_1_pmp_4_cfg_a = io_dpath_pmp_4_cfg_a;
	assign io_requestor_1_pmp_4_cfg_x = io_dpath_pmp_4_cfg_x;
	assign io_requestor_1_pmp_4_cfg_w = io_dpath_pmp_4_cfg_w;
	assign io_requestor_1_pmp_4_cfg_r = io_dpath_pmp_4_cfg_r;
	assign io_requestor_1_pmp_4_addr = io_dpath_pmp_4_addr;
	assign io_requestor_1_pmp_4_mask = io_dpath_pmp_4_mask;
	assign io_requestor_1_pmp_5_cfg_l = io_dpath_pmp_5_cfg_l;
	assign io_requestor_1_pmp_5_cfg_a = io_dpath_pmp_5_cfg_a;
	assign io_requestor_1_pmp_5_cfg_x = io_dpath_pmp_5_cfg_x;
	assign io_requestor_1_pmp_5_cfg_w = io_dpath_pmp_5_cfg_w;
	assign io_requestor_1_pmp_5_cfg_r = io_dpath_pmp_5_cfg_r;
	assign io_requestor_1_pmp_5_addr = io_dpath_pmp_5_addr;
	assign io_requestor_1_pmp_5_mask = io_dpath_pmp_5_mask;
	assign io_requestor_1_pmp_6_cfg_l = io_dpath_pmp_6_cfg_l;
	assign io_requestor_1_pmp_6_cfg_a = io_dpath_pmp_6_cfg_a;
	assign io_requestor_1_pmp_6_cfg_x = io_dpath_pmp_6_cfg_x;
	assign io_requestor_1_pmp_6_cfg_w = io_dpath_pmp_6_cfg_w;
	assign io_requestor_1_pmp_6_cfg_r = io_dpath_pmp_6_cfg_r;
	assign io_requestor_1_pmp_6_addr = io_dpath_pmp_6_addr;
	assign io_requestor_1_pmp_6_mask = io_dpath_pmp_6_mask;
	assign io_requestor_1_pmp_7_cfg_l = io_dpath_pmp_7_cfg_l;
	assign io_requestor_1_pmp_7_cfg_a = io_dpath_pmp_7_cfg_a;
	assign io_requestor_1_pmp_7_cfg_x = io_dpath_pmp_7_cfg_x;
	assign io_requestor_1_pmp_7_cfg_w = io_dpath_pmp_7_cfg_w;
	assign io_requestor_1_pmp_7_cfg_r = io_dpath_pmp_7_cfg_r;
	assign io_requestor_1_pmp_7_addr = io_dpath_pmp_7_addr;
	assign io_requestor_1_pmp_7_mask = io_dpath_pmp_7_mask;
	assign io_requestor_1_customCSRs_csrs_0_value = io_dpath_customCSRs_csrs_0_value;
	assign io_dpath_perf_l2hit = 1'h0;
	assign io_dpath_perf_pte_miss = 1'h0;
	assign io_dpath_perf_pte_hit = 1'h0;
	assign l2_tlb_ram_RW0_clk = clock;
	assign l2_tlb_ram_RW0_wdata_0 = {_T_133, _T_132};
	assign state_barrier_io_x = (3'h0 == state ? state : _GEN_2207);
	assign r_pte_barrier_io_x_ppn = ((state == 3'h7) & _T_199 ? pte_2_ppn : r_pte_ppn);
	assign r_pte_barrier_io_x_d = r_pte_d;
	assign r_pte_barrier_io_x_a = r_pte_a;
	assign r_pte_barrier_io_x_u = r_pte_u;
	assign r_pte_barrier_io_x_x = r_pte_x;
	assign r_pte_barrier_io_x_w = r_pte_w;
	assign r_pte_barrier_io_x_r = r_pte_r;
	always @(posedge clock) begin
		if (reset)
			state <= 3'h0;
		else
			state <= state_barrier_io_y;
		r_pte_ppn <= r_pte_barrier_io_y_ppn;
		r_pte_d <= r_pte_barrier_io_y_d;
		r_pte_a <= r_pte_barrier_io_y_a;
		r_pte_u <= r_pte_barrier_io_y_u;
		r_pte_x <= r_pte_barrier_io_y_x;
		r_pte_w <= r_pte_barrier_io_y_w;
		r_pte_r <= r_pte_barrier_io_y_r;
	end
endmodule
module RVCExpander (
	io_in,
	io_out_bits,
	io_out_rd,
	io_out_rs1,
	io_out_rs2,
	io_rvc
);
	input [31:0] io_in;
	output wire [31:0] io_out_bits;
	output wire [4:0] io_out_rd;
	output wire [4:0] io_out_rs1;
	output wire [4:0] io_out_rs2;
	output wire io_rvc;
	wire [6:0] io_out_s_opc = (|io_in[12:5] ? 7'h13 : 7'h1f);
	wire [4:0] _io_out_s_T_6 = {2'h1, io_in[4:2]};
	wire [29:0] _io_out_s_T_7 = {io_in[10:7], io_in[12:11], io_in[5], io_in[6], 2'h0, 5'h02, 3'h0, 2'h1, io_in[4:2], io_out_s_opc};
	wire [7:0] _io_out_s_T_15 = {io_in[6:5], io_in[12:10], 3'h0};
	wire [4:0] _io_out_s_T_17 = {2'h1, io_in[9:7]};
	wire [27:0] _io_out_s_T_20 = {io_in[6:5], io_in[12:10], 3'h0, 2'h1, io_in[9:7], 3'h3, 2'h1, io_in[4:2], 7'h07};
	wire [6:0] _io_out_s_T_31 = {io_in[5], io_in[12:10], io_in[6], 2'h0};
	wire [26:0] _io_out_s_T_36 = {io_in[5], io_in[12:10], io_in[6], 2'h0, 2'h1, io_in[9:7], 3'h2, 2'h1, io_in[4:2], 7'h03};
	wire [26:0] _io_out_s_T_52 = {io_in[5], io_in[12:10], io_in[6], 2'h0, 2'h1, io_in[9:7], 3'h2, 2'h1, io_in[4:2], 7'h07};
	wire [26:0] _io_out_s_T_74 = {_io_out_s_T_31[6:5], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, _io_out_s_T_31[4:0], 7'h3f};
	wire [27:0] _io_out_s_T_94 = {_io_out_s_T_15[7:5], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h3, _io_out_s_T_15[4:0], 7'h27};
	wire [26:0] _io_out_s_T_116 = {_io_out_s_T_31[6:5], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, _io_out_s_T_31[4:0], 7'h23};
	wire [26:0] _io_out_s_T_138 = {_io_out_s_T_31[6:5], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, _io_out_s_T_31[4:0], 7'h27};
	wire [6:0] _io_out_s_T_148 = (io_in[12] ? 7'h7f : 7'h00);
	wire [11:0] _io_out_s_T_150 = {_io_out_s_T_148, io_in[6:2]};
	wire [31:0] io_out_s_8_bits = {_io_out_s_T_148, io_in[6:2], io_in[11:7], 3'h0, io_in[11:7], 7'h13};
	wire [9:0] _io_out_s_T_161 = (io_in[12] ? 10'h3ff : 10'h000);
	wire [20:0] _io_out_s_T_169 = {_io_out_s_T_161, io_in[8], io_in[10:9], io_in[6], io_in[7], io_in[2], io_in[11], io_in[5:3], 1'h0};
	wire [31:0] io_out_s_9_bits = {_io_out_s_T_169[20], _io_out_s_T_169[10:1], _io_out_s_T_169[11], _io_out_s_T_169[19:12], 5'h01, 7'h6f};
	wire [31:0] io_out_s_10_bits = {_io_out_s_T_148, io_in[6:2], 5'h00, 3'h0, io_in[11:7], 7'h13};
	wire _io_out_s_opc_T_7 = |_io_out_s_T_150;
	wire [6:0] io_out_s_opc_1 = (|_io_out_s_T_150 ? 7'h37 : 7'h3f);
	wire [14:0] _io_out_s_me_T_2 = (io_in[12] ? 15'h7fff : 15'h0000);
	wire [31:0] _io_out_s_me_T_4 = {_io_out_s_me_T_2, io_in[6:2], 12'h000};
	wire [31:0] io_out_s_me_bits = {_io_out_s_me_T_4[31:12], io_in[11:7], io_out_s_opc_1};
	wire [6:0] io_out_s_opc_2 = (_io_out_s_opc_T_7 ? 7'h13 : 7'h1f);
	wire [2:0] _io_out_s_T_230 = (io_in[12] ? 3'h7 : 3'h0);
	wire [31:0] io_out_s_res_bits = {_io_out_s_T_230, io_in[4:3], io_in[5], io_in[2], io_in[6], 4'h0, io_in[11:7], 3'h0, io_in[11:7], io_out_s_opc_2};
	wire [31:0] io_out_s_11_bits = ((io_in[11:7] == 5'h00) | (io_in[11:7] == 5'h02) ? io_out_s_res_bits : io_out_s_me_bits);
	wire [4:0] io_out_s_11_rd = ((io_in[11:7] == 5'h00) | (io_in[11:7] == 5'h02) ? io_in[11:7] : io_in[11:7]);
	wire [4:0] io_out_s_11_rs2 = ((io_in[11:7] == 5'h00) | (io_in[11:7] == 5'h02) ? _io_out_s_T_6 : _io_out_s_T_6);
	wire [25:0] _io_out_s_T_251 = {io_in[12], io_in[6:2], 2'h1, io_in[9:7], 3'h5, 2'h1, io_in[9:7], 7'h13};
	wire [30:0] _GEN_0 = {5'd0, _io_out_s_T_251};
	wire [30:0] _io_out_s_T_260 = _GEN_0 | 31'h40000000;
	wire [31:0] _io_out_s_T_270 = {_io_out_s_T_148, io_in[6:2], 2'h1, io_in[9:7], 3'h7, 2'h1, io_in[9:7], 7'h13};
	wire [2:0] _io_out_s_funct_T_2 = {io_in[12], io_in[6:5]};
	wire [2:0] _io_out_s_funct_T_4 = (_io_out_s_funct_T_2 == 3'h1 ? 3'h4 : 3'h0);
	wire [2:0] _io_out_s_funct_T_6 = (_io_out_s_funct_T_2 == 3'h2 ? 3'h6 : _io_out_s_funct_T_4);
	wire [2:0] _io_out_s_funct_T_8 = (_io_out_s_funct_T_2 == 3'h3 ? 3'h7 : _io_out_s_funct_T_6);
	wire [2:0] _io_out_s_funct_T_10 = (_io_out_s_funct_T_2 == 3'h4 ? 3'h0 : _io_out_s_funct_T_8);
	wire [2:0] _io_out_s_funct_T_12 = (_io_out_s_funct_T_2 == 3'h5 ? 3'h0 : _io_out_s_funct_T_10);
	wire [2:0] _io_out_s_funct_T_14 = (_io_out_s_funct_T_2 == 3'h6 ? 3'h2 : _io_out_s_funct_T_12);
	wire [2:0] io_out_s_funct = (_io_out_s_funct_T_2 == 3'h7 ? 3'h3 : _io_out_s_funct_T_14);
	wire [30:0] io_out_s_sub = (io_in[6:5] == 2'h0 ? 31'h40000000 : 31'h00000000);
	wire [6:0] io_out_s_opc_3 = (io_in[12] ? 7'h3b : 7'h33);
	wire [24:0] _io_out_s_T_277 = {2'h1, io_in[4:2], 2'h1, io_in[9:7], io_out_s_funct, 2'h1, io_in[9:7], io_out_s_opc_3};
	wire [30:0] _GEN_1 = {6'd0, _io_out_s_T_277};
	wire [30:0] _io_out_s_T_278 = _GEN_1 | io_out_s_sub;
	wire [30:0] _io_out_s_T_281 = (io_in[11:10] == 2'h1 ? _io_out_s_T_260 : {5'd0, _io_out_s_T_251});
	wire [31:0] _io_out_s_T_283 = (io_in[11:10] == 2'h2 ? _io_out_s_T_270 : {1'd0, _io_out_s_T_281});
	wire [31:0] io_out_s_12_bits = (io_in[11:10] == 2'h3 ? {1'd0, _io_out_s_T_278} : _io_out_s_T_283);
	wire [31:0] io_out_s_13_bits = {_io_out_s_T_169[20], _io_out_s_T_169[10:1], _io_out_s_T_169[11], _io_out_s_T_169[19:12], 5'h00, 7'h6f};
	wire [4:0] _io_out_s_T_349 = (io_in[12] ? 5'h1f : 5'h00);
	wire [12:0] _io_out_s_T_354 = {_io_out_s_T_349, io_in[6:5], io_in[2], io_in[11:10], io_in[4:3], 1'h0};
	wire [31:0] io_out_s_14_bits = {_io_out_s_T_354[12], _io_out_s_T_354[10:5], 5'h00, 2'h1, io_in[9:7], 3'h0, _io_out_s_T_354[4:1], _io_out_s_T_354[11], 7'h63};
	wire [31:0] io_out_s_15_bits = {_io_out_s_T_354[12], _io_out_s_T_354[10:5], 5'h00, 2'h1, io_in[9:7], 3'h1, _io_out_s_T_354[4:1], _io_out_s_T_354[11], 7'h63};
	wire _io_out_s_load_opc_T_1 = |io_in[11:7];
	wire [6:0] io_out_s_load_opc = (|io_in[11:7] ? 7'h03 : 7'h1f);
	wire [25:0] _io_out_s_T_438 = {io_in[12], io_in[6:2], io_in[11:7], 3'h1, io_in[11:7], 7'h13};
	wire [28:0] _io_out_s_T_448 = {io_in[4:2], io_in[12], io_in[6:5], 3'h0, 5'h02, 3'h3, io_in[11:7], 7'h07};
	wire [27:0] _io_out_s_T_457 = {io_in[3:2], io_in[12], io_in[6:4], 2'h0, 5'h02, 3'h2, io_in[11:7], io_out_s_load_opc};
	wire [27:0] _io_out_s_T_466 = {io_in[3:2], io_in[12], io_in[6:4], 2'h0, 5'h02, 3'h2, io_in[11:7], 7'h07};
	wire [24:0] _io_out_s_mv_T_2 = {io_in[6:2], 5'h00, 3'h0, io_in[11:7], 7'h33};
	wire [24:0] _io_out_s_add_T_3 = {io_in[6:2], io_in[11:7], 3'h0, io_in[11:7], 7'h33};
	wire [24:0] io_out_s_jr = {io_in[6:2], io_in[11:7], 3'h0, 12'h067};
	wire [24:0] io_out_s_reserved = {io_out_s_jr[24:7], 7'h1f};
	wire [24:0] _io_out_s_jr_reserved_T_2 = (_io_out_s_load_opc_T_1 ? io_out_s_jr : io_out_s_reserved);
	wire _io_out_s_jr_mv_T_1 = |io_in[6:2];
	wire [31:0] io_out_s_mv_bits = {7'd0, _io_out_s_mv_T_2};
	wire [31:0] io_out_s_jr_reserved_bits = {7'd0, _io_out_s_jr_reserved_T_2};
	wire [31:0] io_out_s_jr_mv_bits = (|io_in[6:2] ? io_out_s_mv_bits : io_out_s_jr_reserved_bits);
	wire [4:0] io_out_s_jr_mv_rd = (|io_in[6:2] ? io_in[11:7] : 5'h00);
	wire [4:0] io_out_s_jr_mv_rs1 = (|io_in[6:2] ? 5'h00 : io_in[11:7]);
	wire [4:0] io_out_s_jr_mv_rs2 = (|io_in[6:2] ? io_in[6:2] : io_in[6:2]);
	wire [24:0] io_out_s_jalr = {io_in[6:2], io_in[11:7], 3'h0, 12'h0e7};
	wire [24:0] _io_out_s_ebreak_T_1 = {io_out_s_jr[24:7], 7'h73};
	wire [24:0] io_out_s_ebreak = _io_out_s_ebreak_T_1 | 25'h0100000;
	wire [24:0] _io_out_s_jalr_ebreak_T_2 = (_io_out_s_load_opc_T_1 ? io_out_s_jalr : io_out_s_ebreak);
	wire [31:0] io_out_s_add_bits = {7'd0, _io_out_s_add_T_3};
	wire [31:0] io_out_s_jalr_ebreak_bits = {7'd0, _io_out_s_jalr_ebreak_T_2};
	wire [31:0] io_out_s_jalr_add_bits = (_io_out_s_jr_mv_T_1 ? io_out_s_add_bits : io_out_s_jalr_ebreak_bits);
	wire [4:0] io_out_s_jalr_add_rd = (_io_out_s_jr_mv_T_1 ? io_in[11:7] : 5'h01);
	wire [4:0] io_out_s_jalr_add_rs1 = (_io_out_s_jr_mv_T_1 ? io_in[11:7] : io_in[11:7]);
	wire [31:0] io_out_s_20_bits = (io_in[12] ? io_out_s_jalr_add_bits : io_out_s_jr_mv_bits);
	wire [4:0] io_out_s_20_rd = (io_in[12] ? io_out_s_jalr_add_rd : io_out_s_jr_mv_rd);
	wire [4:0] io_out_s_20_rs1 = (io_in[12] ? io_out_s_jalr_add_rs1 : io_out_s_jr_mv_rs1);
	wire [4:0] io_out_s_20_rs2 = (io_in[12] ? io_out_s_jr_mv_rs2 : io_out_s_jr_mv_rs2);
	wire [8:0] _io_out_s_T_473 = {io_in[9:7], io_in[12:10], 3'h0};
	wire [28:0] _io_out_s_T_480 = {_io_out_s_T_473[8:5], io_in[6:2], 5'h02, 3'h3, _io_out_s_T_473[4:0], 7'h27};
	wire [7:0] _io_out_s_T_486 = {io_in[8:7], io_in[12:9], 2'h0};
	wire [27:0] _io_out_s_T_493 = {_io_out_s_T_486[7:5], io_in[6:2], 5'h02, 3'h2, _io_out_s_T_486[4:0], 7'h23};
	wire [27:0] _io_out_s_T_506 = {_io_out_s_T_486[7:5], io_in[6:2], 5'h02, 3'h2, _io_out_s_T_486[4:0], 7'h27};
	wire [4:0] io_out_s_24_rs1 = io_in[19:15];
	wire [4:0] io_out_s_24_rs2 = io_in[24:20];
	wire [4:0] _io_out_T_2 = {io_in[1:0], io_in[15:13]};
	wire [31:0] io_out_s_1_bits = {4'd0, _io_out_s_T_20};
	wire [31:0] io_out_s_0_bits = {2'd0, _io_out_s_T_7};
	wire [31:0] _io_out_T_4_bits = (_io_out_T_2 == 5'h01 ? io_out_s_1_bits : io_out_s_0_bits);
	wire [4:0] _io_out_T_4_rd = (_io_out_T_2 == 5'h01 ? _io_out_s_T_6 : _io_out_s_T_6);
	wire [4:0] _io_out_T_4_rs1 = (_io_out_T_2 == 5'h01 ? _io_out_s_T_17 : 5'h02);
	wire [31:0] io_out_s_2_bits = {5'd0, _io_out_s_T_36};
	wire [31:0] _io_out_T_6_bits = (_io_out_T_2 == 5'h02 ? io_out_s_2_bits : _io_out_T_4_bits);
	wire [4:0] _io_out_T_6_rd = (_io_out_T_2 == 5'h02 ? _io_out_s_T_6 : _io_out_T_4_rd);
	wire [4:0] _io_out_T_6_rs1 = (_io_out_T_2 == 5'h02 ? _io_out_s_T_17 : _io_out_T_4_rs1);
	wire [31:0] io_out_s_3_bits = {5'd0, _io_out_s_T_52};
	wire [31:0] _io_out_T_8_bits = (_io_out_T_2 == 5'h03 ? io_out_s_3_bits : _io_out_T_6_bits);
	wire [4:0] _io_out_T_8_rd = (_io_out_T_2 == 5'h03 ? _io_out_s_T_6 : _io_out_T_6_rd);
	wire [4:0] _io_out_T_8_rs1 = (_io_out_T_2 == 5'h03 ? _io_out_s_T_17 : _io_out_T_6_rs1);
	wire [31:0] io_out_s_4_bits = {5'd0, _io_out_s_T_74};
	wire [31:0] _io_out_T_10_bits = (_io_out_T_2 == 5'h04 ? io_out_s_4_bits : _io_out_T_8_bits);
	wire [4:0] _io_out_T_10_rd = (_io_out_T_2 == 5'h04 ? _io_out_s_T_6 : _io_out_T_8_rd);
	wire [4:0] _io_out_T_10_rs1 = (_io_out_T_2 == 5'h04 ? _io_out_s_T_17 : _io_out_T_8_rs1);
	wire [31:0] io_out_s_5_bits = {4'd0, _io_out_s_T_94};
	wire [31:0] _io_out_T_12_bits = (_io_out_T_2 == 5'h05 ? io_out_s_5_bits : _io_out_T_10_bits);
	wire [4:0] _io_out_T_12_rd = (_io_out_T_2 == 5'h05 ? _io_out_s_T_6 : _io_out_T_10_rd);
	wire [4:0] _io_out_T_12_rs1 = (_io_out_T_2 == 5'h05 ? _io_out_s_T_17 : _io_out_T_10_rs1);
	wire [31:0] io_out_s_6_bits = {5'd0, _io_out_s_T_116};
	wire [31:0] _io_out_T_14_bits = (_io_out_T_2 == 5'h06 ? io_out_s_6_bits : _io_out_T_12_bits);
	wire [4:0] _io_out_T_14_rd = (_io_out_T_2 == 5'h06 ? _io_out_s_T_6 : _io_out_T_12_rd);
	wire [4:0] _io_out_T_14_rs1 = (_io_out_T_2 == 5'h06 ? _io_out_s_T_17 : _io_out_T_12_rs1);
	wire [31:0] io_out_s_7_bits = {5'd0, _io_out_s_T_138};
	wire [31:0] _io_out_T_16_bits = (_io_out_T_2 == 5'h07 ? io_out_s_7_bits : _io_out_T_14_bits);
	wire [4:0] _io_out_T_16_rd = (_io_out_T_2 == 5'h07 ? _io_out_s_T_6 : _io_out_T_14_rd);
	wire [4:0] _io_out_T_16_rs1 = (_io_out_T_2 == 5'h07 ? _io_out_s_T_17 : _io_out_T_14_rs1);
	wire [31:0] _io_out_T_18_bits = (_io_out_T_2 == 5'h08 ? io_out_s_8_bits : _io_out_T_16_bits);
	wire [4:0] _io_out_T_18_rd = (_io_out_T_2 == 5'h08 ? io_in[11:7] : _io_out_T_16_rd);
	wire [4:0] _io_out_T_18_rs1 = (_io_out_T_2 == 5'h08 ? io_in[11:7] : _io_out_T_16_rs1);
	wire [4:0] _io_out_T_18_rs2 = (_io_out_T_2 == 5'h08 ? _io_out_s_T_6 : _io_out_T_16_rd);
	wire [31:0] _io_out_T_20_bits = (_io_out_T_2 == 5'h09 ? io_out_s_9_bits : _io_out_T_18_bits);
	wire [4:0] _io_out_T_20_rd = (_io_out_T_2 == 5'h09 ? 5'h01 : _io_out_T_18_rd);
	wire [4:0] _io_out_T_20_rs1 = (_io_out_T_2 == 5'h09 ? io_in[11:7] : _io_out_T_18_rs1);
	wire [4:0] _io_out_T_20_rs2 = (_io_out_T_2 == 5'h09 ? _io_out_s_T_6 : _io_out_T_18_rs2);
	wire [31:0] _io_out_T_22_bits = (_io_out_T_2 == 5'h0a ? io_out_s_10_bits : _io_out_T_20_bits);
	wire [4:0] _io_out_T_22_rd = (_io_out_T_2 == 5'h0a ? io_in[11:7] : _io_out_T_20_rd);
	wire [4:0] _io_out_T_22_rs1 = (_io_out_T_2 == 5'h0a ? 5'h00 : _io_out_T_20_rs1);
	wire [4:0] _io_out_T_22_rs2 = (_io_out_T_2 == 5'h0a ? _io_out_s_T_6 : _io_out_T_20_rs2);
	wire [31:0] _io_out_T_24_bits = (_io_out_T_2 == 5'h0b ? io_out_s_11_bits : _io_out_T_22_bits);
	wire [4:0] _io_out_T_24_rd = (_io_out_T_2 == 5'h0b ? io_out_s_11_rd : _io_out_T_22_rd);
	wire [4:0] _io_out_T_24_rs1 = (_io_out_T_2 == 5'h0b ? io_out_s_11_rd : _io_out_T_22_rs1);
	wire [4:0] _io_out_T_24_rs2 = (_io_out_T_2 == 5'h0b ? io_out_s_11_rs2 : _io_out_T_22_rs2);
	wire [31:0] _io_out_T_26_bits = (_io_out_T_2 == 5'h0c ? io_out_s_12_bits : _io_out_T_24_bits);
	wire [4:0] _io_out_T_26_rd = (_io_out_T_2 == 5'h0c ? _io_out_s_T_17 : _io_out_T_24_rd);
	wire [4:0] _io_out_T_26_rs1 = (_io_out_T_2 == 5'h0c ? _io_out_s_T_17 : _io_out_T_24_rs1);
	wire [4:0] _io_out_T_26_rs2 = (_io_out_T_2 == 5'h0c ? _io_out_s_T_6 : _io_out_T_24_rs2);
	wire [31:0] _io_out_T_28_bits = (_io_out_T_2 == 5'h0d ? io_out_s_13_bits : _io_out_T_26_bits);
	wire [4:0] _io_out_T_28_rd = (_io_out_T_2 == 5'h0d ? 5'h00 : _io_out_T_26_rd);
	wire [4:0] _io_out_T_28_rs1 = (_io_out_T_2 == 5'h0d ? _io_out_s_T_17 : _io_out_T_26_rs1);
	wire [4:0] _io_out_T_28_rs2 = (_io_out_T_2 == 5'h0d ? _io_out_s_T_6 : _io_out_T_26_rs2);
	wire [31:0] _io_out_T_30_bits = (_io_out_T_2 == 5'h0e ? io_out_s_14_bits : _io_out_T_28_bits);
	wire [4:0] _io_out_T_30_rd = (_io_out_T_2 == 5'h0e ? _io_out_s_T_17 : _io_out_T_28_rd);
	wire [4:0] _io_out_T_30_rs1 = (_io_out_T_2 == 5'h0e ? _io_out_s_T_17 : _io_out_T_28_rs1);
	wire [4:0] _io_out_T_30_rs2 = (_io_out_T_2 == 5'h0e ? 5'h00 : _io_out_T_28_rs2);
	wire [31:0] _io_out_T_32_bits = (_io_out_T_2 == 5'h0f ? io_out_s_15_bits : _io_out_T_30_bits);
	wire [4:0] _io_out_T_32_rd = (_io_out_T_2 == 5'h0f ? 5'h00 : _io_out_T_30_rd);
	wire [4:0] _io_out_T_32_rs1 = (_io_out_T_2 == 5'h0f ? _io_out_s_T_17 : _io_out_T_30_rs1);
	wire [4:0] _io_out_T_32_rs2 = (_io_out_T_2 == 5'h0f ? 5'h00 : _io_out_T_30_rs2);
	wire [31:0] io_out_s_16_bits = {6'd0, _io_out_s_T_438};
	wire [31:0] _io_out_T_34_bits = (_io_out_T_2 == 5'h10 ? io_out_s_16_bits : _io_out_T_32_bits);
	wire [4:0] _io_out_T_34_rd = (_io_out_T_2 == 5'h10 ? io_in[11:7] : _io_out_T_32_rd);
	wire [4:0] _io_out_T_34_rs1 = (_io_out_T_2 == 5'h10 ? io_in[11:7] : _io_out_T_32_rs1);
	wire [4:0] _io_out_T_34_rs2 = (_io_out_T_2 == 5'h10 ? io_in[6:2] : _io_out_T_32_rs2);
	wire [31:0] io_out_s_17_bits = {3'd0, _io_out_s_T_448};
	wire [31:0] _io_out_T_36_bits = (_io_out_T_2 == 5'h11 ? io_out_s_17_bits : _io_out_T_34_bits);
	wire [4:0] _io_out_T_36_rd = (_io_out_T_2 == 5'h11 ? io_in[11:7] : _io_out_T_34_rd);
	wire [4:0] _io_out_T_36_rs1 = (_io_out_T_2 == 5'h11 ? 5'h02 : _io_out_T_34_rs1);
	wire [4:0] _io_out_T_36_rs2 = (_io_out_T_2 == 5'h11 ? io_in[6:2] : _io_out_T_34_rs2);
	wire [31:0] io_out_s_18_bits = {4'd0, _io_out_s_T_457};
	wire [31:0] _io_out_T_38_bits = (_io_out_T_2 == 5'h12 ? io_out_s_18_bits : _io_out_T_36_bits);
	wire [4:0] _io_out_T_38_rd = (_io_out_T_2 == 5'h12 ? io_in[11:7] : _io_out_T_36_rd);
	wire [4:0] _io_out_T_38_rs1 = (_io_out_T_2 == 5'h12 ? 5'h02 : _io_out_T_36_rs1);
	wire [4:0] _io_out_T_38_rs2 = (_io_out_T_2 == 5'h12 ? io_in[6:2] : _io_out_T_36_rs2);
	wire [31:0] io_out_s_19_bits = {4'd0, _io_out_s_T_466};
	wire [31:0] _io_out_T_40_bits = (_io_out_T_2 == 5'h13 ? io_out_s_19_bits : _io_out_T_38_bits);
	wire [4:0] _io_out_T_40_rd = (_io_out_T_2 == 5'h13 ? io_in[11:7] : _io_out_T_38_rd);
	wire [4:0] _io_out_T_40_rs1 = (_io_out_T_2 == 5'h13 ? 5'h02 : _io_out_T_38_rs1);
	wire [4:0] _io_out_T_40_rs2 = (_io_out_T_2 == 5'h13 ? io_in[6:2] : _io_out_T_38_rs2);
	wire [31:0] _io_out_T_42_bits = (_io_out_T_2 == 5'h14 ? io_out_s_20_bits : _io_out_T_40_bits);
	wire [4:0] _io_out_T_42_rd = (_io_out_T_2 == 5'h14 ? io_out_s_20_rd : _io_out_T_40_rd);
	wire [4:0] _io_out_T_42_rs1 = (_io_out_T_2 == 5'h14 ? io_out_s_20_rs1 : _io_out_T_40_rs1);
	wire [4:0] _io_out_T_42_rs2 = (_io_out_T_2 == 5'h14 ? io_out_s_20_rs2 : _io_out_T_40_rs2);
	wire [31:0] io_out_s_21_bits = {3'd0, _io_out_s_T_480};
	wire [31:0] _io_out_T_44_bits = (_io_out_T_2 == 5'h15 ? io_out_s_21_bits : _io_out_T_42_bits);
	wire [4:0] _io_out_T_44_rd = (_io_out_T_2 == 5'h15 ? io_in[11:7] : _io_out_T_42_rd);
	wire [4:0] _io_out_T_44_rs1 = (_io_out_T_2 == 5'h15 ? 5'h02 : _io_out_T_42_rs1);
	wire [4:0] _io_out_T_44_rs2 = (_io_out_T_2 == 5'h15 ? io_in[6:2] : _io_out_T_42_rs2);
	wire [31:0] io_out_s_22_bits = {4'd0, _io_out_s_T_493};
	wire [31:0] _io_out_T_46_bits = (_io_out_T_2 == 5'h16 ? io_out_s_22_bits : _io_out_T_44_bits);
	wire [4:0] _io_out_T_46_rd = (_io_out_T_2 == 5'h16 ? io_in[11:7] : _io_out_T_44_rd);
	wire [4:0] _io_out_T_46_rs1 = (_io_out_T_2 == 5'h16 ? 5'h02 : _io_out_T_44_rs1);
	wire [4:0] _io_out_T_46_rs2 = (_io_out_T_2 == 5'h16 ? io_in[6:2] : _io_out_T_44_rs2);
	wire [31:0] io_out_s_23_bits = {4'd0, _io_out_s_T_506};
	wire [31:0] _io_out_T_48_bits = (_io_out_T_2 == 5'h17 ? io_out_s_23_bits : _io_out_T_46_bits);
	wire [4:0] _io_out_T_48_rd = (_io_out_T_2 == 5'h17 ? io_in[11:7] : _io_out_T_46_rd);
	wire [4:0] _io_out_T_48_rs1 = (_io_out_T_2 == 5'h17 ? 5'h02 : _io_out_T_46_rs1);
	wire [4:0] _io_out_T_48_rs2 = (_io_out_T_2 == 5'h17 ? io_in[6:2] : _io_out_T_46_rs2);
	wire [31:0] _io_out_T_50_bits = (_io_out_T_2 == 5'h18 ? io_in : _io_out_T_48_bits);
	wire [4:0] _io_out_T_50_rd = (_io_out_T_2 == 5'h18 ? io_in[11:7] : _io_out_T_48_rd);
	wire [4:0] _io_out_T_50_rs1 = (_io_out_T_2 == 5'h18 ? io_out_s_24_rs1 : _io_out_T_48_rs1);
	wire [4:0] _io_out_T_50_rs2 = (_io_out_T_2 == 5'h18 ? io_out_s_24_rs2 : _io_out_T_48_rs2);
	wire [31:0] _io_out_T_52_bits = (_io_out_T_2 == 5'h19 ? io_in : _io_out_T_50_bits);
	wire [4:0] _io_out_T_52_rd = (_io_out_T_2 == 5'h19 ? io_in[11:7] : _io_out_T_50_rd);
	wire [4:0] _io_out_T_52_rs1 = (_io_out_T_2 == 5'h19 ? io_out_s_24_rs1 : _io_out_T_50_rs1);
	wire [4:0] _io_out_T_52_rs2 = (_io_out_T_2 == 5'h19 ? io_out_s_24_rs2 : _io_out_T_50_rs2);
	wire [31:0] _io_out_T_54_bits = (_io_out_T_2 == 5'h1a ? io_in : _io_out_T_52_bits);
	wire [4:0] _io_out_T_54_rd = (_io_out_T_2 == 5'h1a ? io_in[11:7] : _io_out_T_52_rd);
	wire [4:0] _io_out_T_54_rs1 = (_io_out_T_2 == 5'h1a ? io_out_s_24_rs1 : _io_out_T_52_rs1);
	wire [4:0] _io_out_T_54_rs2 = (_io_out_T_2 == 5'h1a ? io_out_s_24_rs2 : _io_out_T_52_rs2);
	wire [31:0] _io_out_T_56_bits = (_io_out_T_2 == 5'h1b ? io_in : _io_out_T_54_bits);
	wire [4:0] _io_out_T_56_rd = (_io_out_T_2 == 5'h1b ? io_in[11:7] : _io_out_T_54_rd);
	wire [4:0] _io_out_T_56_rs1 = (_io_out_T_2 == 5'h1b ? io_out_s_24_rs1 : _io_out_T_54_rs1);
	wire [4:0] _io_out_T_56_rs2 = (_io_out_T_2 == 5'h1b ? io_out_s_24_rs2 : _io_out_T_54_rs2);
	wire [31:0] _io_out_T_58_bits = (_io_out_T_2 == 5'h1c ? io_in : _io_out_T_56_bits);
	wire [4:0] _io_out_T_58_rd = (_io_out_T_2 == 5'h1c ? io_in[11:7] : _io_out_T_56_rd);
	wire [4:0] _io_out_T_58_rs1 = (_io_out_T_2 == 5'h1c ? io_out_s_24_rs1 : _io_out_T_56_rs1);
	wire [4:0] _io_out_T_58_rs2 = (_io_out_T_2 == 5'h1c ? io_out_s_24_rs2 : _io_out_T_56_rs2);
	wire [31:0] _io_out_T_60_bits = (_io_out_T_2 == 5'h1d ? io_in : _io_out_T_58_bits);
	wire [4:0] _io_out_T_60_rd = (_io_out_T_2 == 5'h1d ? io_in[11:7] : _io_out_T_58_rd);
	wire [4:0] _io_out_T_60_rs1 = (_io_out_T_2 == 5'h1d ? io_out_s_24_rs1 : _io_out_T_58_rs1);
	wire [4:0] _io_out_T_60_rs2 = (_io_out_T_2 == 5'h1d ? io_out_s_24_rs2 : _io_out_T_58_rs2);
	wire [31:0] _io_out_T_62_bits = (_io_out_T_2 == 5'h1e ? io_in : _io_out_T_60_bits);
	wire [4:0] _io_out_T_62_rd = (_io_out_T_2 == 5'h1e ? io_in[11:7] : _io_out_T_60_rd);
	wire [4:0] _io_out_T_62_rs1 = (_io_out_T_2 == 5'h1e ? io_out_s_24_rs1 : _io_out_T_60_rs1);
	wire [4:0] _io_out_T_62_rs2 = (_io_out_T_2 == 5'h1e ? io_out_s_24_rs2 : _io_out_T_60_rs2);
	assign io_out_bits = (_io_out_T_2 == 5'h1f ? io_in : _io_out_T_62_bits);
	assign io_out_rd = (_io_out_T_2 == 5'h1f ? io_in[11:7] : _io_out_T_62_rd);
	assign io_out_rs1 = (_io_out_T_2 == 5'h1f ? io_out_s_24_rs1 : _io_out_T_62_rs1);
	assign io_out_rs2 = (_io_out_T_2 == 5'h1f ? io_out_s_24_rs2 : _io_out_T_62_rs2);
	assign io_rvc = io_in[1:0] != 2'h3;
endmodule
module IBuf (
	clock,
	reset,
	io_imem_ready,
	io_imem_valid,
	io_imem_bits_pc,
	io_imem_bits_data,
	io_imem_bits_xcpt_ae_inst,
	io_imem_bits_replay,
	io_kill,
	io_pc,
	io_inst_0_ready,
	io_inst_0_valid,
	io_inst_0_bits_xcpt0_ae_inst,
	io_inst_0_bits_xcpt1_pf_inst,
	io_inst_0_bits_xcpt1_gf_inst,
	io_inst_0_bits_xcpt1_ae_inst,
	io_inst_0_bits_replay,
	io_inst_0_bits_rvc,
	io_inst_0_bits_inst_bits,
	io_inst_0_bits_inst_rd,
	io_inst_0_bits_inst_rs1,
	io_inst_0_bits_inst_rs2,
	io_inst_0_bits_raw
);
	input clock;
	input reset;
	output wire io_imem_ready;
	input io_imem_valid;
	input [31:0] io_imem_bits_pc;
	input [31:0] io_imem_bits_data;
	input io_imem_bits_xcpt_ae_inst;
	input io_imem_bits_replay;
	input io_kill;
	output wire [31:0] io_pc;
	input io_inst_0_ready;
	output wire io_inst_0_valid;
	output wire io_inst_0_bits_xcpt0_ae_inst;
	output wire io_inst_0_bits_xcpt1_pf_inst;
	output wire io_inst_0_bits_xcpt1_gf_inst;
	output wire io_inst_0_bits_xcpt1_ae_inst;
	output wire io_inst_0_bits_replay;
	output wire io_inst_0_bits_rvc;
	output wire [31:0] io_inst_0_bits_inst_bits;
	output wire [4:0] io_inst_0_bits_inst_rd;
	output wire [4:0] io_inst_0_bits_inst_rs1;
	output wire [4:0] io_inst_0_bits_inst_rs2;
	output wire [31:0] io_inst_0_bits_raw;
	wire [31:0] exp_io_in;
	wire [31:0] exp_io_out_bits;
	wire [4:0] exp_io_out_rd;
	wire [4:0] exp_io_out_rs1;
	wire [4:0] exp_io_out_rs2;
	wire exp_io_rvc;
	reg nBufValid;
	reg [31:0] buf__pc;
	reg [31:0] buf__data;
	reg buf__xcpt_ae_inst;
	reg buf__replay;
	wire pcWordBits = io_imem_bits_pc[1];
	wire [1:0] _GEN_58 = {1'd0, pcWordBits};
	wire [1:0] nIC = 2'h2 - _GEN_58;
	wire [1:0] _nValid_T = (io_imem_valid ? nIC : 2'h0);
	wire [1:0] _GEN_59 = {1'd0, nBufValid};
	wire [1:0] nValid = _nValid_T + _GEN_59;
	wire [3:0] _valid_T = 4'h1 << nValid;
	wire [3:0] _valid_T_2 = _valid_T - 4'h1;
	wire [1:0] valid = _valid_T_2[1:0];
	wire [1:0] _full_insn_T_2 = {1'd0, valid[1]};
	wire [1:0] _bufMask_T = 2'h1 << nBufValid;
	wire [1:0] bufMask = _bufMask_T - 2'h1;
	wire [1:0] buf_replay = (buf__replay ? bufMask : 2'h0);
	wire full_insn = (exp_io_rvc | _full_insn_T_2[0]) | buf_replay[0];
	wire [1:0] _nReady_T_4 = (exp_io_rvc ? 2'h1 : 2'h2);
	wire [1:0] nReady = (full_insn ? _nReady_T_4 : 2'h0);
	wire [1:0] nICReady = nReady - _GEN_59;
	wire _io_imem_ready_T = nReady >= _GEN_59;
	wire [1:0] _io_imem_ready_T_4 = nIC - nICReady;
	wire _io_imem_ready_T_5 = 2'h1 >= _io_imem_ready_T_4;
	wire _nBufValid_T_2 = _io_imem_ready_T | ~nBufValid;
	wire [1:0] _nBufValid_T_4 = _GEN_59 - nReady;
	wire [1:0] _nBufValid_T_5 = (_nBufValid_T_2 ? 2'h0 : _nBufValid_T_4);
	wire [1:0] shamt = _GEN_58 + nICReady;
	wire [63:0] buf_data_data = {io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data};
	wire [5:0] _buf_data_T = {shamt, 4'h0};
	wire [63:0] _buf_data_T_1 = buf_data_data >> _buf_data_T;
	wire [31:0] _buf_pc_T_1 = io_imem_bits_pc & 32'hfffffffc;
	wire [2:0] _buf_pc_T_2 = {nICReady, 1'h0};
	wire [31:0] _GEN_67 = {29'd0, _buf_pc_T_2};
	wire [31:0] _buf_pc_T_4 = io_imem_bits_pc + _GEN_67;
	wire [31:0] _buf_pc_T_5 = _buf_pc_T_4 & 32'h00000003;
	wire [31:0] _buf_pc_T_6 = _buf_pc_T_1 | _buf_pc_T_5;
	wire [1:0] _GEN_0 = (((io_imem_valid & _io_imem_ready_T) & (nICReady < nIC)) & _io_imem_ready_T_5 ? _io_imem_ready_T_4 : _nBufValid_T_5);
	wire [1:0] _GEN_24 = (io_inst_0_ready ? _GEN_0 : {1'd0, nBufValid});
	wire [1:0] _GEN_48 = (io_kill ? 2'h0 : _GEN_24);
	wire [1:0] _icShiftAmt_T_1 = 2'h2 + _GEN_59;
	wire [1:0] icShiftAmt = _icShiftAmt_T_1 - _GEN_58;
	wire [63:0] _icData_T_2 = {io_imem_bits_data, io_imem_bits_data[15:0], io_imem_bits_data[15:0]};
	wire [127:0] icData_data = {_icData_T_2[63:48], _icData_T_2[63:48], _icData_T_2[63:48], _icData_T_2[63:48], io_imem_bits_data, io_imem_bits_data[15:0], io_imem_bits_data[15:0]};
	wire [5:0] _icData_T_3 = {icShiftAmt, 4'h0};
	wire [190:0] _GEN_1 = {63'd0, icData_data};
	wire [190:0] _icData_T_4 = _GEN_1 << _icData_T_3;
	wire [31:0] icData = _icData_T_4[95:64];
	wire [4:0] _icMask_T_1 = {nBufValid, 4'h0};
	wire [62:0] _icMask_T_2 = 63'h00000000ffffffff << _icMask_T_1;
	wire [31:0] icMask = _icMask_T_2[31:0];
	wire [31:0] _inst_T = icData & icMask;
	wire [31:0] _inst_T_1 = ~icMask;
	wire [31:0] _inst_T_2 = buf__data & _inst_T_1;
	wire xcpt_1_ae_inst = (bufMask[1] ? buf__xcpt_ae_inst : io_imem_bits_xcpt_ae_inst);
	wire [1:0] _ic_replay_T = ~bufMask;
	wire [1:0] _ic_replay_T_1 = valid & _ic_replay_T;
	wire [1:0] _ic_replay_T_2 = (io_imem_bits_replay ? _ic_replay_T_1 : 2'h0);
	wire [1:0] ic_replay = buf_replay | _ic_replay_T_2;
	wire [1:0] _replay_T_5 = {1'd0, ic_replay[1]};
	wire [2:0] _io_inst_0_bits_xcpt1_T_4 = {2'h0, xcpt_1_ae_inst};
	wire [2:0] _io_inst_0_bits_xcpt1_T_5 = (exp_io_rvc ? 3'h0 : _io_inst_0_bits_xcpt1_T_4);
	RVCExpander exp(
		.io_in(exp_io_in),
		.io_out_bits(exp_io_out_bits),
		.io_out_rd(exp_io_out_rd),
		.io_out_rs1(exp_io_out_rs1),
		.io_out_rs2(exp_io_out_rs2),
		.io_rvc(exp_io_rvc)
	);
	assign io_imem_ready = (io_inst_0_ready & (nReady >= _GEN_59)) & ((nICReady >= nIC) | (2'h1 >= _io_imem_ready_T_4));
	assign io_pc = (nBufValid > 1'h0 ? buf__pc : io_imem_bits_pc);
	assign io_inst_0_valid = valid[0] & full_insn;
	assign io_inst_0_bits_xcpt0_ae_inst = (bufMask[0] ? buf__xcpt_ae_inst : io_imem_bits_xcpt_ae_inst);
	assign io_inst_0_bits_xcpt1_pf_inst = _io_inst_0_bits_xcpt1_T_5[2];
	assign io_inst_0_bits_xcpt1_gf_inst = _io_inst_0_bits_xcpt1_T_5[1];
	assign io_inst_0_bits_xcpt1_ae_inst = _io_inst_0_bits_xcpt1_T_5[0];
	assign io_inst_0_bits_replay = ic_replay[0] | (~exp_io_rvc & _replay_T_5[0]);
	assign io_inst_0_bits_rvc = exp_io_rvc;
	assign io_inst_0_bits_inst_bits = exp_io_out_bits;
	assign io_inst_0_bits_inst_rd = exp_io_out_rd;
	assign io_inst_0_bits_inst_rs1 = exp_io_out_rs1;
	assign io_inst_0_bits_inst_rs2 = exp_io_out_rs2;
	assign io_inst_0_bits_raw = _inst_T | _inst_T_2;
	assign exp_io_in = _inst_T | _inst_T_2;
	always @(posedge clock) begin
		if (reset)
			nBufValid <= 1'h0;
		else
			nBufValid <= _GEN_48[0];
		if (io_inst_0_ready)
			if (((io_imem_valid & _io_imem_ready_T) & (nICReady < nIC)) & _io_imem_ready_T_5)
				buf__pc <= _buf_pc_T_6;
		if (io_inst_0_ready)
			if (((io_imem_valid & _io_imem_ready_T) & (nICReady < nIC)) & _io_imem_ready_T_5)
				buf__data <= {16'd0, _buf_data_T_1[15:0]};
		if (io_inst_0_ready)
			if (((io_imem_valid & _io_imem_ready_T) & (nICReady < nIC)) & _io_imem_ready_T_5)
				buf__xcpt_ae_inst <= io_imem_bits_xcpt_ae_inst;
		if (io_inst_0_ready)
			if (((io_imem_valid & _io_imem_ready_T) & (nICReady < nIC)) & _io_imem_ready_T_5)
				buf__replay <= io_imem_bits_replay;
	end
endmodule
module CSRFile (
	clock,
	reset,
	io_ungated_clock,
	io_interrupts_debug,
	io_interrupts_mtip,
	io_interrupts_msip,
	io_interrupts_meip,
	io_hartid,
	io_rw_addr,
	io_rw_cmd,
	io_rw_rdata,
	io_rw_wdata,
	io_decode_0_inst,
	io_decode_0_fp_illegal,
	io_decode_0_fp_csr,
	io_decode_0_read_illegal,
	io_decode_0_write_illegal,
	io_decode_0_write_flush,
	io_decode_0_system_illegal,
	io_csr_stall,
	io_eret,
	io_singleStep,
	io_status_debug,
	io_status_cease,
	io_status_wfi,
	io_status_isa,
	io_status_dprv,
	io_status_dv,
	io_status_prv,
	io_status_v,
	io_status_sd,
	io_status_zero2,
	io_status_mpv,
	io_status_gva,
	io_status_mbe,
	io_status_sbe,
	io_status_sxl,
	io_status_uxl,
	io_status_sd_rv32,
	io_status_zero1,
	io_status_tsr,
	io_status_tw,
	io_status_tvm,
	io_status_mxr,
	io_status_sum,
	io_status_mprv,
	io_status_xs,
	io_status_fs,
	io_status_mpp,
	io_status_vs,
	io_status_spp,
	io_status_mpie,
	io_status_ube,
	io_status_spie,
	io_status_upie,
	io_status_mie,
	io_status_hie,
	io_status_sie,
	io_status_uie,
	io_evec,
	io_exception,
	io_retire,
	io_cause,
	io_pc,
	io_tval,
	io_gva,
	io_time,
	io_interrupt,
	io_interrupt_cause,
	io_bp_0_control_action,
	io_bp_0_control_tmatch,
	io_bp_0_control_x,
	io_bp_0_control_w,
	io_bp_0_control_r,
	io_bp_0_address,
	io_pmp_0_cfg_l,
	io_pmp_0_cfg_a,
	io_pmp_0_cfg_x,
	io_pmp_0_cfg_w,
	io_pmp_0_cfg_r,
	io_pmp_0_addr,
	io_pmp_0_mask,
	io_pmp_1_cfg_l,
	io_pmp_1_cfg_a,
	io_pmp_1_cfg_x,
	io_pmp_1_cfg_w,
	io_pmp_1_cfg_r,
	io_pmp_1_addr,
	io_pmp_1_mask,
	io_pmp_2_cfg_l,
	io_pmp_2_cfg_a,
	io_pmp_2_cfg_x,
	io_pmp_2_cfg_w,
	io_pmp_2_cfg_r,
	io_pmp_2_addr,
	io_pmp_2_mask,
	io_pmp_3_cfg_l,
	io_pmp_3_cfg_a,
	io_pmp_3_cfg_x,
	io_pmp_3_cfg_w,
	io_pmp_3_cfg_r,
	io_pmp_3_addr,
	io_pmp_3_mask,
	io_pmp_4_cfg_l,
	io_pmp_4_cfg_a,
	io_pmp_4_cfg_x,
	io_pmp_4_cfg_w,
	io_pmp_4_cfg_r,
	io_pmp_4_addr,
	io_pmp_4_mask,
	io_pmp_5_cfg_l,
	io_pmp_5_cfg_a,
	io_pmp_5_cfg_x,
	io_pmp_5_cfg_w,
	io_pmp_5_cfg_r,
	io_pmp_5_addr,
	io_pmp_5_mask,
	io_pmp_6_cfg_l,
	io_pmp_6_cfg_a,
	io_pmp_6_cfg_x,
	io_pmp_6_cfg_w,
	io_pmp_6_cfg_r,
	io_pmp_6_addr,
	io_pmp_6_mask,
	io_pmp_7_cfg_l,
	io_pmp_7_cfg_a,
	io_pmp_7_cfg_x,
	io_pmp_7_cfg_w,
	io_pmp_7_cfg_r,
	io_pmp_7_addr,
	io_pmp_7_mask,
	io_inhibit_cycle,
	io_inst_0,
	io_trace_0_valid,
	io_trace_0_iaddr,
	io_trace_0_insn,
	io_trace_0_exception,
	io_customCSRs_0_value
);
	input clock;
	input reset;
	input io_ungated_clock;
	input io_interrupts_debug;
	input io_interrupts_mtip;
	input io_interrupts_msip;
	input io_interrupts_meip;
	input io_hartid;
	input [11:0] io_rw_addr;
	input [2:0] io_rw_cmd;
	output wire [31:0] io_rw_rdata;
	input [31:0] io_rw_wdata;
	input [31:0] io_decode_0_inst;
	output wire io_decode_0_fp_illegal;
	output wire io_decode_0_fp_csr;
	output wire io_decode_0_read_illegal;
	output wire io_decode_0_write_illegal;
	output wire io_decode_0_write_flush;
	output wire io_decode_0_system_illegal;
	output wire io_csr_stall;
	output wire io_eret;
	output wire io_singleStep;
	output wire io_status_debug;
	output wire io_status_cease;
	output wire io_status_wfi;
	output wire [31:0] io_status_isa;
	output wire [1:0] io_status_dprv;
	output wire io_status_dv;
	output wire [1:0] io_status_prv;
	output wire io_status_v;
	output wire io_status_sd;
	output wire [22:0] io_status_zero2;
	output wire io_status_mpv;
	output wire io_status_gva;
	output wire io_status_mbe;
	output wire io_status_sbe;
	output wire [1:0] io_status_sxl;
	output wire [1:0] io_status_uxl;
	output wire io_status_sd_rv32;
	output wire [7:0] io_status_zero1;
	output wire io_status_tsr;
	output wire io_status_tw;
	output wire io_status_tvm;
	output wire io_status_mxr;
	output wire io_status_sum;
	output wire io_status_mprv;
	output wire [1:0] io_status_xs;
	output wire [1:0] io_status_fs;
	output wire [1:0] io_status_mpp;
	output wire [1:0] io_status_vs;
	output wire io_status_spp;
	output wire io_status_mpie;
	output wire io_status_ube;
	output wire io_status_spie;
	output wire io_status_upie;
	output wire io_status_mie;
	output wire io_status_hie;
	output wire io_status_sie;
	output wire io_status_uie;
	output wire [31:0] io_evec;
	input io_exception;
	input io_retire;
	input [31:0] io_cause;
	input [31:0] io_pc;
	input [31:0] io_tval;
	input io_gva;
	output wire [31:0] io_time;
	output wire io_interrupt;
	output wire [31:0] io_interrupt_cause;
	output wire io_bp_0_control_action;
	output wire [1:0] io_bp_0_control_tmatch;
	output wire io_bp_0_control_x;
	output wire io_bp_0_control_w;
	output wire io_bp_0_control_r;
	output wire [31:0] io_bp_0_address;
	output wire io_pmp_0_cfg_l;
	output wire [1:0] io_pmp_0_cfg_a;
	output wire io_pmp_0_cfg_x;
	output wire io_pmp_0_cfg_w;
	output wire io_pmp_0_cfg_r;
	output wire [29:0] io_pmp_0_addr;
	output wire [31:0] io_pmp_0_mask;
	output wire io_pmp_1_cfg_l;
	output wire [1:0] io_pmp_1_cfg_a;
	output wire io_pmp_1_cfg_x;
	output wire io_pmp_1_cfg_w;
	output wire io_pmp_1_cfg_r;
	output wire [29:0] io_pmp_1_addr;
	output wire [31:0] io_pmp_1_mask;
	output wire io_pmp_2_cfg_l;
	output wire [1:0] io_pmp_2_cfg_a;
	output wire io_pmp_2_cfg_x;
	output wire io_pmp_2_cfg_w;
	output wire io_pmp_2_cfg_r;
	output wire [29:0] io_pmp_2_addr;
	output wire [31:0] io_pmp_2_mask;
	output wire io_pmp_3_cfg_l;
	output wire [1:0] io_pmp_3_cfg_a;
	output wire io_pmp_3_cfg_x;
	output wire io_pmp_3_cfg_w;
	output wire io_pmp_3_cfg_r;
	output wire [29:0] io_pmp_3_addr;
	output wire [31:0] io_pmp_3_mask;
	output wire io_pmp_4_cfg_l;
	output wire [1:0] io_pmp_4_cfg_a;
	output wire io_pmp_4_cfg_x;
	output wire io_pmp_4_cfg_w;
	output wire io_pmp_4_cfg_r;
	output wire [29:0] io_pmp_4_addr;
	output wire [31:0] io_pmp_4_mask;
	output wire io_pmp_5_cfg_l;
	output wire [1:0] io_pmp_5_cfg_a;
	output wire io_pmp_5_cfg_x;
	output wire io_pmp_5_cfg_w;
	output wire io_pmp_5_cfg_r;
	output wire [29:0] io_pmp_5_addr;
	output wire [31:0] io_pmp_5_mask;
	output wire io_pmp_6_cfg_l;
	output wire [1:0] io_pmp_6_cfg_a;
	output wire io_pmp_6_cfg_x;
	output wire io_pmp_6_cfg_w;
	output wire io_pmp_6_cfg_r;
	output wire [29:0] io_pmp_6_addr;
	output wire [31:0] io_pmp_6_mask;
	output wire io_pmp_7_cfg_l;
	output wire [1:0] io_pmp_7_cfg_a;
	output wire io_pmp_7_cfg_x;
	output wire io_pmp_7_cfg_w;
	output wire io_pmp_7_cfg_r;
	output wire [29:0] io_pmp_7_addr;
	output wire [31:0] io_pmp_7_mask;
	output wire io_inhibit_cycle;
	input [31:0] io_inst_0;
	output wire io_trace_0_valid;
	output wire [31:0] io_trace_0_iaddr;
	output wire [31:0] io_trace_0_insn;
	output wire io_trace_0_exception;
	output wire [31:0] io_customCSRs_0_value;
	reg reg_mstatus_gva;
	reg reg_mstatus_spp;
	reg reg_mstatus_mpie;
	reg reg_mstatus_mie;
	reg reg_dcsr_ebreakm;
	reg [2:0] reg_dcsr_cause;
	reg reg_dcsr_step;
	reg reg_debug;
	reg [31:0] reg_dpc;
	reg [31:0] reg_dscratch;
	reg reg_singleStepped;
	reg reg_bp_0_control_dmode;
	reg reg_bp_0_control_action;
	reg [1:0] reg_bp_0_control_tmatch;
	reg reg_bp_0_control_x;
	reg reg_bp_0_control_w;
	reg reg_bp_0_control_r;
	reg [31:0] reg_bp_0_address;
	reg reg_pmp_0_cfg_l;
	reg [1:0] reg_pmp_0_cfg_a;
	reg reg_pmp_0_cfg_x;
	reg reg_pmp_0_cfg_w;
	reg reg_pmp_0_cfg_r;
	reg [29:0] reg_pmp_0_addr;
	reg reg_pmp_1_cfg_l;
	reg [1:0] reg_pmp_1_cfg_a;
	reg reg_pmp_1_cfg_x;
	reg reg_pmp_1_cfg_w;
	reg reg_pmp_1_cfg_r;
	reg [29:0] reg_pmp_1_addr;
	reg reg_pmp_2_cfg_l;
	reg [1:0] reg_pmp_2_cfg_a;
	reg reg_pmp_2_cfg_x;
	reg reg_pmp_2_cfg_w;
	reg reg_pmp_2_cfg_r;
	reg [29:0] reg_pmp_2_addr;
	reg reg_pmp_3_cfg_l;
	reg [1:0] reg_pmp_3_cfg_a;
	reg reg_pmp_3_cfg_x;
	reg reg_pmp_3_cfg_w;
	reg reg_pmp_3_cfg_r;
	reg [29:0] reg_pmp_3_addr;
	reg reg_pmp_4_cfg_l;
	reg [1:0] reg_pmp_4_cfg_a;
	reg reg_pmp_4_cfg_x;
	reg reg_pmp_4_cfg_w;
	reg reg_pmp_4_cfg_r;
	reg [29:0] reg_pmp_4_addr;
	reg reg_pmp_5_cfg_l;
	reg [1:0] reg_pmp_5_cfg_a;
	reg reg_pmp_5_cfg_x;
	reg reg_pmp_5_cfg_w;
	reg reg_pmp_5_cfg_r;
	reg [29:0] reg_pmp_5_addr;
	reg reg_pmp_6_cfg_l;
	reg [1:0] reg_pmp_6_cfg_a;
	reg reg_pmp_6_cfg_x;
	reg reg_pmp_6_cfg_w;
	reg reg_pmp_6_cfg_r;
	reg [29:0] reg_pmp_6_addr;
	reg reg_pmp_7_cfg_l;
	reg [1:0] reg_pmp_7_cfg_a;
	reg reg_pmp_7_cfg_x;
	reg reg_pmp_7_cfg_w;
	reg reg_pmp_7_cfg_r;
	reg [29:0] reg_pmp_7_addr;
	reg [31:0] reg_mie;
	reg [31:0] reg_mepc;
	reg [31:0] reg_mcause;
	reg [31:0] reg_mtval;
	reg [31:0] reg_mscratch;
	reg [31:0] reg_mtvec;
	reg reg_wfi;
	reg [2:0] reg_mcountinhibit;
	wire x79 = reg_mcountinhibit[2];
	reg [5:0] small_;
	wire [5:0] _GEN_34 = {5'd0, io_retire};
	wire [6:0] nextSmall = small_ + _GEN_34;
	wire _T_14 = ~x79;
	wire [6:0] _GEN_0 = (~x79 ? nextSmall : {1'd0, small_});
	reg [57:0] large_;
	wire [57:0] _large_r_T_1 = large_ + 58'h000000000000001;
	wire [57:0] _GEN_1 = (nextSmall[6] & _T_14 ? _large_r_T_1 : large_);
	wire [63:0] value = {large_, small_};
	wire x86 = ~io_csr_stall;
	reg [5:0] small_1;
	wire [5:0] _GEN_35 = {5'd0, x86};
	wire [6:0] nextSmall_1 = small_1 + _GEN_35;
	wire _T_15 = ~reg_mcountinhibit[0];
	wire [6:0] _GEN_2 = (~reg_mcountinhibit[0] ? nextSmall_1 : {1'd0, small_1});
	reg [57:0] large_1;
	wire [57:0] _large_r_T_3 = large_1 + 58'h000000000000001;
	wire [57:0] _GEN_3 = (nextSmall_1[6] & _T_15 ? _large_r_T_3 : large_1);
	wire [63:0] value_1 = {large_1, small_1};
	wire [15:0] _read_mip_T = {4'h0, io_interrupts_meip, 1'h0, 2'h0, io_interrupts_mtip, 1'h0, 2'h0, io_interrupts_msip, 1'h0, 2'h0};
	wire [15:0] read_mip = _read_mip_T & 16'h0888;
	wire [31:0] _GEN_40 = {16'd0, read_mip};
	wire [31:0] pending_interrupts = _GEN_40 & reg_mie;
	wire [14:0] d_interrupts = {io_interrupts_debug, 14'h0000};
	wire [31:0] _m_interrupts_T_3 = ~pending_interrupts;
	wire [31:0] _m_interrupts_T_5 = ~_m_interrupts_T_3;
	wire [31:0] m_interrupts = (reg_mstatus_mie ? _m_interrupts_T_5 : 32'h00000000);
	wire _any_T_78 = ((((((((((((((d_interrupts[14] | d_interrupts[13]) | d_interrupts[12]) | d_interrupts[11]) | d_interrupts[3]) | d_interrupts[7]) | d_interrupts[9]) | d_interrupts[1]) | d_interrupts[5]) | d_interrupts[10]) | d_interrupts[2]) | d_interrupts[6]) | d_interrupts[8]) | d_interrupts[0]) | d_interrupts[4]) | m_interrupts[15];
	wire anyInterrupt = ((((((((((((((_any_T_78 | m_interrupts[14]) | m_interrupts[13]) | m_interrupts[12]) | m_interrupts[11]) | m_interrupts[3]) | m_interrupts[7]) | m_interrupts[9]) | m_interrupts[1]) | m_interrupts[5]) | m_interrupts[10]) | m_interrupts[2]) | m_interrupts[6]) | m_interrupts[8]) | m_interrupts[0]) | m_interrupts[4];
	wire [3:0] _which_T_95 = (m_interrupts[0] ? 4'h0 : 4'h4);
	wire [3:0] _which_T_96 = (m_interrupts[8] ? 4'h8 : _which_T_95);
	wire [3:0] _which_T_97 = (m_interrupts[6] ? 4'h6 : _which_T_96);
	wire [3:0] _which_T_98 = (m_interrupts[2] ? 4'h2 : _which_T_97);
	wire [3:0] _which_T_99 = (m_interrupts[10] ? 4'ha : _which_T_98);
	wire [3:0] _which_T_100 = (m_interrupts[5] ? 4'h5 : _which_T_99);
	wire [3:0] _which_T_101 = (m_interrupts[1] ? 4'h1 : _which_T_100);
	wire [3:0] _which_T_102 = (m_interrupts[9] ? 4'h9 : _which_T_101);
	wire [3:0] _which_T_103 = (m_interrupts[7] ? 4'h7 : _which_T_102);
	wire [3:0] _which_T_104 = (m_interrupts[3] ? 4'h3 : _which_T_103);
	wire [3:0] _which_T_105 = (m_interrupts[11] ? 4'hb : _which_T_104);
	wire [3:0] _which_T_106 = (m_interrupts[12] ? 4'hc : _which_T_105);
	wire [3:0] _which_T_107 = (m_interrupts[13] ? 4'hd : _which_T_106);
	wire [3:0] _which_T_108 = (m_interrupts[14] ? 4'he : _which_T_107);
	wire [3:0] _which_T_109 = (m_interrupts[15] ? 4'hf : _which_T_108);
	wire [3:0] _which_T_111 = (d_interrupts[4] ? 4'h4 : _which_T_109);
	wire [3:0] _which_T_112 = (d_interrupts[0] ? 4'h0 : _which_T_111);
	wire [3:0] _which_T_113 = (d_interrupts[8] ? 4'h8 : _which_T_112);
	wire [3:0] _which_T_114 = (d_interrupts[6] ? 4'h6 : _which_T_113);
	wire [3:0] _which_T_115 = (d_interrupts[2] ? 4'h2 : _which_T_114);
	wire [3:0] _which_T_116 = (d_interrupts[10] ? 4'ha : _which_T_115);
	wire [3:0] _which_T_117 = (d_interrupts[5] ? 4'h5 : _which_T_116);
	wire [3:0] _which_T_118 = (d_interrupts[1] ? 4'h1 : _which_T_117);
	wire [3:0] _which_T_119 = (d_interrupts[9] ? 4'h9 : _which_T_118);
	wire [3:0] _which_T_120 = (d_interrupts[7] ? 4'h7 : _which_T_119);
	wire [3:0] _which_T_121 = (d_interrupts[3] ? 4'h3 : _which_T_120);
	wire [3:0] _which_T_122 = (d_interrupts[11] ? 4'hb : _which_T_121);
	wire [3:0] _which_T_123 = (d_interrupts[12] ? 4'hc : _which_T_122);
	wire [3:0] _which_T_124 = (d_interrupts[13] ? 4'hd : _which_T_123);
	wire [3:0] whichInterrupt = (d_interrupts[14] ? 4'he : _which_T_124);
	wire [31:0] _GEN_41 = {28'd0, whichInterrupt};
	wire _io_interrupt_T = ~io_singleStep;
	wire [30:0] pmp_mask_base = {reg_pmp_0_addr, reg_pmp_0_cfg_a[0]};
	wire [30:0] _pmp_mask_T_1 = pmp_mask_base + 31'h00000001;
	wire [30:0] _pmp_mask_T_2 = ~_pmp_mask_T_1;
	wire [30:0] _pmp_mask_T_3 = pmp_mask_base & _pmp_mask_T_2;
	wire [32:0] _pmp_mask_T_4 = {_pmp_mask_T_3, 2'h3};
	wire [30:0] pmp_mask_base_1 = {reg_pmp_1_addr, reg_pmp_1_cfg_a[0]};
	wire [30:0] _pmp_mask_T_6 = pmp_mask_base_1 + 31'h00000001;
	wire [30:0] _pmp_mask_T_7 = ~_pmp_mask_T_6;
	wire [30:0] _pmp_mask_T_8 = pmp_mask_base_1 & _pmp_mask_T_7;
	wire [32:0] _pmp_mask_T_9 = {_pmp_mask_T_8, 2'h3};
	wire [30:0] pmp_mask_base_2 = {reg_pmp_2_addr, reg_pmp_2_cfg_a[0]};
	wire [30:0] _pmp_mask_T_11 = pmp_mask_base_2 + 31'h00000001;
	wire [30:0] _pmp_mask_T_12 = ~_pmp_mask_T_11;
	wire [30:0] _pmp_mask_T_13 = pmp_mask_base_2 & _pmp_mask_T_12;
	wire [32:0] _pmp_mask_T_14 = {_pmp_mask_T_13, 2'h3};
	wire [30:0] pmp_mask_base_3 = {reg_pmp_3_addr, reg_pmp_3_cfg_a[0]};
	wire [30:0] _pmp_mask_T_16 = pmp_mask_base_3 + 31'h00000001;
	wire [30:0] _pmp_mask_T_17 = ~_pmp_mask_T_16;
	wire [30:0] _pmp_mask_T_18 = pmp_mask_base_3 & _pmp_mask_T_17;
	wire [32:0] _pmp_mask_T_19 = {_pmp_mask_T_18, 2'h3};
	wire [30:0] pmp_mask_base_4 = {reg_pmp_4_addr, reg_pmp_4_cfg_a[0]};
	wire [30:0] _pmp_mask_T_21 = pmp_mask_base_4 + 31'h00000001;
	wire [30:0] _pmp_mask_T_22 = ~_pmp_mask_T_21;
	wire [30:0] _pmp_mask_T_23 = pmp_mask_base_4 & _pmp_mask_T_22;
	wire [32:0] _pmp_mask_T_24 = {_pmp_mask_T_23, 2'h3};
	wire [30:0] pmp_mask_base_5 = {reg_pmp_5_addr, reg_pmp_5_cfg_a[0]};
	wire [30:0] _pmp_mask_T_26 = pmp_mask_base_5 + 31'h00000001;
	wire [30:0] _pmp_mask_T_27 = ~_pmp_mask_T_26;
	wire [30:0] _pmp_mask_T_28 = pmp_mask_base_5 & _pmp_mask_T_27;
	wire [32:0] _pmp_mask_T_29 = {_pmp_mask_T_28, 2'h3};
	wire [30:0] pmp_mask_base_6 = {reg_pmp_6_addr, reg_pmp_6_cfg_a[0]};
	wire [30:0] _pmp_mask_T_31 = pmp_mask_base_6 + 31'h00000001;
	wire [30:0] _pmp_mask_T_32 = ~_pmp_mask_T_31;
	wire [30:0] _pmp_mask_T_33 = pmp_mask_base_6 & _pmp_mask_T_32;
	wire [32:0] _pmp_mask_T_34 = {_pmp_mask_T_33, 2'h3};
	wire [30:0] pmp_mask_base_7 = {reg_pmp_7_addr, reg_pmp_7_cfg_a[0]};
	wire [30:0] _pmp_mask_T_36 = pmp_mask_base_7 + 31'h00000001;
	wire [30:0] _pmp_mask_T_37 = ~_pmp_mask_T_36;
	wire [30:0] _pmp_mask_T_38 = pmp_mask_base_7 & _pmp_mask_T_37;
	wire [32:0] _pmp_mask_T_39 = {_pmp_mask_T_38, 2'h3};
	reg [31:0] reg_misa;
	wire [8:0] read_mstatus_lo_lo = {io_status_spp, io_status_mpie, io_status_ube, io_status_spie, io_status_upie, io_status_mie, io_status_hie, io_status_sie, io_status_uie};
	wire [21:0] read_mstatus_lo = {io_status_tw, io_status_tvm, io_status_mxr, io_status_sum, io_status_mprv, io_status_xs, io_status_fs, io_status_mpp, io_status_vs, read_mstatus_lo_lo};
	wire [64:0] read_mstatus_hi_hi = {io_status_debug, io_status_cease, io_status_wfi, io_status_isa, io_status_dprv, io_status_dv, io_status_prv, io_status_v, io_status_sd, io_status_zero2};
	wire [82:0] read_mstatus_hi = {read_mstatus_hi_hi, io_status_mpv, io_status_gva, io_status_mbe, io_status_sbe, io_status_sxl, io_status_uxl, io_status_sd_rv32, io_status_zero1, io_status_tsr};
	wire [104:0] _read_mstatus_T = {read_mstatus_hi, read_mstatus_lo};
	wire [31:0] read_mstatus = _read_mstatus_T[31:0];
	wire [6:0] _read_mtvec_T_1 = (reg_mtvec[0] ? 7'h7e : 7'h02);
	wire [31:0] _read_mtvec_T_3 = {25'd0, _read_mtvec_T_1};
	wire [31:0] _read_mtvec_T_4 = ~_read_mtvec_T_3;
	wire [31:0] read_mtvec = reg_mtvec & _read_mtvec_T_4;
	wire [6:0] lo_4 = {4'h8, reg_bp_0_control_x, reg_bp_0_control_w, reg_bp_0_control_r};
	wire [31:0] _T_16 = {4'h2, reg_bp_0_control_dmode, 14'h0400, reg_bp_0_control_action, 1'h0, 2'h0, reg_bp_0_control_tmatch, lo_4};
	wire [31:0] _T_18 = ~reg_mepc;
	wire [1:0] _T_20 = (reg_misa[2] ? 2'h1 : 2'h3);
	wire [31:0] _GEN_586 = {30'd0, _T_20};
	wire [31:0] _T_21 = _T_18 | _GEN_586;
	wire [31:0] _T_22 = ~_T_21;
	wire [31:0] _T_23 = {16'h4000, reg_dcsr_ebreakm, 4'h0, 2'h0, reg_dcsr_cause, 1'h0, 2'h0, reg_dcsr_step, 2'h3};
	wire [31:0] _T_24 = ~reg_dpc;
	wire [31:0] _T_27 = _T_24 | _GEN_586;
	wire [31:0] _T_28 = ~_T_27;
	wire [7:0] _T_60 = {reg_pmp_0_cfg_l, 2'h0, reg_pmp_0_cfg_a, reg_pmp_0_cfg_x, reg_pmp_0_cfg_w, reg_pmp_0_cfg_r};
	wire [7:0] _T_62 = {reg_pmp_2_cfg_l, 2'h0, reg_pmp_2_cfg_a, reg_pmp_2_cfg_x, reg_pmp_2_cfg_w, reg_pmp_2_cfg_r};
	wire [15:0] lo_11 = {reg_pmp_1_cfg_l, 2'h0, reg_pmp_1_cfg_a, reg_pmp_1_cfg_x, reg_pmp_1_cfg_w, reg_pmp_1_cfg_r, _T_60};
	wire [31:0] _T_64 = {reg_pmp_3_cfg_l, 2'h0, reg_pmp_3_cfg_a, reg_pmp_3_cfg_x, reg_pmp_3_cfg_w, reg_pmp_3_cfg_r, _T_62, lo_11};
	wire [7:0] _T_65 = {reg_pmp_4_cfg_l, 2'h0, reg_pmp_4_cfg_a, reg_pmp_4_cfg_x, reg_pmp_4_cfg_w, reg_pmp_4_cfg_r};
	wire [7:0] _T_67 = {reg_pmp_6_cfg_l, 2'h0, reg_pmp_6_cfg_a, reg_pmp_6_cfg_x, reg_pmp_6_cfg_w, reg_pmp_6_cfg_r};
	wire [15:0] lo_16 = {reg_pmp_5_cfg_l, 2'h0, reg_pmp_5_cfg_a, reg_pmp_5_cfg_x, reg_pmp_5_cfg_w, reg_pmp_5_cfg_r, _T_65};
	wire [31:0] _T_69 = {reg_pmp_7_cfg_l, 2'h0, reg_pmp_7_cfg_a, reg_pmp_7_cfg_x, reg_pmp_7_cfg_w, reg_pmp_7_cfg_r, _T_67, lo_16};
	reg [31:0] reg_custom_0;
	wire [12:0] addr = {io_status_v, io_rw_addr};
	wire [12:0] _decoded_T = addr & 13'h0413;
	wire [12:0] _decoded_T_2 = addr & 13'h0453;
	wire decoded_1 = _decoded_T_2 == 13'h0401;
	wire decoded_2 = _decoded_T == 13'h0402;
	wire [12:0] _decoded_T_8 = addr & 13'h0865;
	wire decoded_4 = _decoded_T_8 == 13'h0001;
	wire decoded_5 = _decoded_T_8 == 13'h0000;
	wire [12:0] _decoded_T_12 = addr & 13'h0825;
	wire decoded_6 = _decoded_T_12 == 13'h0005;
	wire [12:0] _decoded_T_14 = addr & 13'h0044;
	wire decoded_7 = _decoded_T_14 == 13'h0044;
	wire decoded_8 = _decoded_T_8 == 13'h0004;
	wire [12:0] _decoded_T_18 = addr & 13'h0047;
	wire decoded_9 = _decoded_T_18 == 13'h0040;
	wire [12:0] _decoded_T_20 = addr & 13'h0443;
	wire decoded_10 = _decoded_T_20 == 13'h0041;
	wire [12:0] _decoded_T_22 = addr & 13'h0823;
	wire decoded_11 = _decoded_T_22 == 13'h0003;
	wire decoded_12 = _decoded_T_22 == 13'h0002;
	wire [12:0] _decoded_T_26 = addr & 13'h0483;
	wire decoded_13 = _decoded_T_26 == 13'h0400;
	wire [12:0] _decoded_T_28 = addr & 13'h0c13;
	wire decoded_14 = _decoded_T_28 == 13'h0410;
	wire [12:0] _decoded_T_30 = addr & 13'h0c11;
	wire decoded_15 = _decoded_T_30 == 13'h0411;
	wire [12:0] _decoded_T_32 = addr & 13'h0c12;
	wire decoded_16 = _decoded_T_32 == 13'h0412;
	wire [12:0] _decoded_T_34 = addr & 13'h00be;
	wire decoded_17 = _decoded_T_34 == 13'h0020;
	wire [12:0] _decoded_T_36 = addr & 13'h089e;
	wire decoded_18 = _decoded_T_36 == 13'h0800;
	wire [12:0] _decoded_T_38 = addr & 13'h00df;
	wire decoded_19 = _decoded_T_38 == 13'h0002;
	wire [12:0] _decoded_T_48 = addr & 13'h089f;
	wire [12:0] _decoded_T_60 = addr & 13'h00bf;
	wire [12:0] _decoded_T_214 = addr & 13'h04be;
	wire decoded_107 = _decoded_T_214 == 13'h0080;
	wire decoded_108 = _decoded_T_60 == 13'h0082;
	wire [12:0] _decoded_T_218 = addr & 13'h0c93;
	wire decoded_109 = _decoded_T_218 == 13'h0080;
	wire decoded_110 = _decoded_T_218 == 13'h0081;
	wire [12:0] _decoded_T_226 = addr & 13'h0c9f;
	wire decoded_113 = _decoded_T_226 == 13'h0090;
	wire decoded_114 = _decoded_T_226 == 13'h0091;
	wire decoded_115 = _decoded_T_226 == 13'h0092;
	wire decoded_116 = _decoded_T_48 == 13'h0093;
	wire [12:0] _decoded_T_234 = addr & 13'h088f;
	wire decoded_117 = _decoded_T_234 == 13'h0084;
	wire decoded_118 = _decoded_T_234 == 13'h0085;
	wire decoded_119 = _decoded_T_234 == 13'h0086;
	wire decoded_120 = _decoded_T_234 == 13'h0087;
	wire [12:0] _decoded_T_258 = addr & 13'h0c20;
	wire decoded_129 = _decoded_T_258 == 13'h0400;
	wire [12:0] _decoded_T_260 = addr & 13'h0485;
	wire decoded_130 = _decoded_T_260 == 13'h0400;
	wire decoded_132 = _decoded_T_26 == 13'h0403;
	wire [31:0] _wdata_T_1 = (io_rw_cmd[1] ? io_rw_rdata : 32'h00000000);
	wire [31:0] _wdata_T_2 = _wdata_T_1 | io_rw_wdata;
	wire [31:0] _wdata_T_5 = (&io_rw_cmd[1:0] ? io_rw_wdata : 32'h00000000);
	wire [31:0] _wdata_T_6 = ~_wdata_T_5;
	wire [31:0] wdata = _wdata_T_2 & _wdata_T_6;
	wire system_insn = io_rw_cmd == 3'h4;
	wire [31:0] _T_213 = {io_rw_addr, 20'h00000};
	wire [31:0] _T_214 = _T_213 & 32'h20100000;
	wire _T_215 = _T_214 == 32'h00000000;
	wire [31:0] _T_217 = _T_213 & 32'h10100000;
	wire _T_218 = _T_217 == 32'h00100000;
	wire [31:0] _T_220 = _T_213 & 32'h20400000;
	wire _T_221 = _T_220 == 32'h20000000;
	wire [31:0] _T_223 = _T_213 & 32'h20200000;
	wire _T_224 = _T_223 == 32'h20000000;
	wire [31:0] _T_226 = _T_213 & 32'h30000000;
	wire _T_227 = _T_226 == 32'h10000000;
	wire insn_call = system_insn & _T_215;
	wire insn_break = system_insn & _T_218;
	wire insn_ret = system_insn & _T_221;
	wire insn_cease = system_insn & _T_224;
	wire insn_wfi = system_insn & _T_227;
	wire [11:0] addr_1 = io_decode_0_inst[31:20];
	wire [31:0] _T_244 = io_decode_0_inst & 32'h20400000;
	wire is_ret = _T_244 == 32'h20000000;
	wire _csr_exists_T_15 = addr_1 == 12'h7b1;
	wire _csr_exists_T_147 = (((((((((((((((addr_1 == 12'h7a0) | (addr_1 == 12'h7a1)) | (addr_1 == 12'h7a2)) | (addr_1 == 12'h7a3)) | (addr_1 == 12'h301)) | (addr_1 == 12'h300)) | (addr_1 == 12'h305)) | (addr_1 == 12'h344)) | (addr_1 == 12'h304)) | (addr_1 == 12'h340)) | (addr_1 == 12'h341)) | (addr_1 == 12'h343)) | (addr_1 == 12'h342)) | (addr_1 == 12'hf14)) | (addr_1 == 12'h7b0)) | _csr_exists_T_15;
	wire _csr_exists_T_162 = ((((((((((((((_csr_exists_T_147 | (addr_1 == 12'h7b2)) | (addr_1 == 12'h320)) | (addr_1 == 12'hb00)) | (addr_1 == 12'hb02)) | (addr_1 == 12'h323)) | (addr_1 == 12'hb03)) | (addr_1 == 12'hb83)) | (addr_1 == 12'h324)) | (addr_1 == 12'hb04)) | (addr_1 == 12'hb84)) | (addr_1 == 12'h325)) | (addr_1 == 12'hb05)) | (addr_1 == 12'hb85)) | (addr_1 == 12'h326)) | (addr_1 == 12'hb06);
	wire _csr_exists_T_177 = ((((((((((((((_csr_exists_T_162 | (addr_1 == 12'hb86)) | (addr_1 == 12'h327)) | (addr_1 == 12'hb07)) | (addr_1 == 12'hb87)) | (addr_1 == 12'h328)) | (addr_1 == 12'hb08)) | (addr_1 == 12'hb88)) | (addr_1 == 12'h329)) | (addr_1 == 12'hb09)) | (addr_1 == 12'hb89)) | (addr_1 == 12'h32a)) | (addr_1 == 12'hb0a)) | (addr_1 == 12'hb8a)) | (addr_1 == 12'h32b)) | (addr_1 == 12'hb0b);
	wire _csr_exists_T_192 = ((((((((((((((_csr_exists_T_177 | (addr_1 == 12'hb8b)) | (addr_1 == 12'h32c)) | (addr_1 == 12'hb0c)) | (addr_1 == 12'hb8c)) | (addr_1 == 12'h32d)) | (addr_1 == 12'hb0d)) | (addr_1 == 12'hb8d)) | (addr_1 == 12'h32e)) | (addr_1 == 12'hb0e)) | (addr_1 == 12'hb8e)) | (addr_1 == 12'h32f)) | (addr_1 == 12'hb0f)) | (addr_1 == 12'hb8f)) | (addr_1 == 12'h330)) | (addr_1 == 12'hb10);
	wire _csr_exists_T_207 = ((((((((((((((_csr_exists_T_192 | (addr_1 == 12'hb90)) | (addr_1 == 12'h331)) | (addr_1 == 12'hb11)) | (addr_1 == 12'hb91)) | (addr_1 == 12'h332)) | (addr_1 == 12'hb12)) | (addr_1 == 12'hb92)) | (addr_1 == 12'h333)) | (addr_1 == 12'hb13)) | (addr_1 == 12'hb93)) | (addr_1 == 12'h334)) | (addr_1 == 12'hb14)) | (addr_1 == 12'hb94)) | (addr_1 == 12'h335)) | (addr_1 == 12'hb15);
	wire _csr_exists_T_222 = ((((((((((((((_csr_exists_T_207 | (addr_1 == 12'hb95)) | (addr_1 == 12'h336)) | (addr_1 == 12'hb16)) | (addr_1 == 12'hb96)) | (addr_1 == 12'h337)) | (addr_1 == 12'hb17)) | (addr_1 == 12'hb97)) | (addr_1 == 12'h338)) | (addr_1 == 12'hb18)) | (addr_1 == 12'hb98)) | (addr_1 == 12'h339)) | (addr_1 == 12'hb19)) | (addr_1 == 12'hb99)) | (addr_1 == 12'h33a)) | (addr_1 == 12'hb1a);
	wire _csr_exists_T_237 = ((((((((((((((_csr_exists_T_222 | (addr_1 == 12'hb9a)) | (addr_1 == 12'h33b)) | (addr_1 == 12'hb1b)) | (addr_1 == 12'hb9b)) | (addr_1 == 12'h33c)) | (addr_1 == 12'hb1c)) | (addr_1 == 12'hb9c)) | (addr_1 == 12'h33d)) | (addr_1 == 12'hb1d)) | (addr_1 == 12'hb9d)) | (addr_1 == 12'h33e)) | (addr_1 == 12'hb1e)) | (addr_1 == 12'hb9e)) | (addr_1 == 12'h33f)) | (addr_1 == 12'hb1f);
	wire _csr_exists_T_252 = ((((((((((((((_csr_exists_T_237 | (addr_1 == 12'hb9f)) | (addr_1 == 12'hb80)) | (addr_1 == 12'hb82)) | (addr_1 == 12'h3a0)) | (addr_1 == 12'h3a1)) | (addr_1 == 12'h3a2)) | (addr_1 == 12'h3a3)) | (addr_1 == 12'h3b0)) | (addr_1 == 12'h3b1)) | (addr_1 == 12'h3b2)) | (addr_1 == 12'h3b3)) | (addr_1 == 12'h3b4)) | (addr_1 == 12'h3b5)) | (addr_1 == 12'h3b6)) | (addr_1 == 12'h3b7);
	wire csr_exists = (((((((((((_csr_exists_T_252 | (addr_1 == 12'h3b8)) | (addr_1 == 12'h3b9)) | (addr_1 == 12'h3ba)) | (addr_1 == 12'h3bb)) | (addr_1 == 12'h3bc)) | (addr_1 == 12'h3bd)) | (addr_1 == 12'h3be)) | (addr_1 == 12'h3bf)) | (addr_1 == 12'h7c1)) | (addr_1 == 12'hf12)) | (addr_1 == 12'hf11)) | (addr_1 == 12'hf13);
	wire _io_decode_0_read_illegal_T_1 = ~csr_exists;
	wire [11:0] _io_decode_0_read_illegal_T_12 = addr_1 & 12'hc10;
	wire _io_decode_0_read_illegal_T_13 = _io_decode_0_read_illegal_T_12 == 12'h410;
	wire _io_decode_0_read_illegal_T_16 = ~reg_debug;
	wire _io_decode_0_read_illegal_T_17 = _io_decode_0_read_illegal_T_13 & ~reg_debug;
	wire _io_decode_0_read_illegal_T_18 = _io_decode_0_read_illegal_T_1 | _io_decode_0_read_illegal_T_17;
	wire _io_decode_0_read_illegal_T_21 = io_decode_0_fp_csr & io_decode_0_fp_illegal;
	wire [11:0] io_decode_0_write_flush_addr_m = addr_1 | 12'h300;
	wire [31:0] _cause_T_5 = (insn_break ? 32'h00000003 : io_cause);
	wire [31:0] cause = (insn_call ? 32'h0000000b : _cause_T_5);
	wire [7:0] cause_lsbs = cause[7:0];
	wire _causeIsDebugInt_T_1 = cause_lsbs == 8'h0e;
	wire causeIsDebugInt = cause[31] & (cause_lsbs == 8'h0e);
	wire _causeIsDebugTrigger_T_1 = ~cause[31];
	wire causeIsDebugTrigger = ~cause[31] & _causeIsDebugInt_T_1;
	wire [3:0] _causeIsDebugBreak_T_3 = {reg_dcsr_ebreakm, 1'h0, 2'h0};
	wire [3:0] _causeIsDebugBreak_T_4 = {3'd0, _causeIsDebugBreak_T_3[3]};
	wire causeIsDebugBreak = (_causeIsDebugTrigger_T_1 & insn_break) & _causeIsDebugBreak_T_4[0];
	wire trapToDebug = (((reg_singleStepped | causeIsDebugInt) | causeIsDebugTrigger) | causeIsDebugBreak) | reg_debug;
	wire [11:0] _debugTVec_T = (insn_break ? 12'h800 : 12'h808);
	wire [11:0] debugTVec = (reg_debug ? _debugTVec_T : 12'h800);
	wire [6:0] notDebugTVec_interruptOffset = {cause[4:0], 2'h0};
	wire [31:0] notDebugTVec_interruptVec = {read_mtvec[31:7], notDebugTVec_interruptOffset};
	wire notDebugTVec_doVector = (read_mtvec[0] & cause[31]) & (cause_lsbs[7:5] == 3'h0);
	wire [31:0] _notDebugTVec_T_1 = {read_mtvec[31:2], 2'h0};
	wire [31:0] notDebugTVec = (notDebugTVec_doVector ? notDebugTVec_interruptVec : _notDebugTVec_T_1);
	wire [31:0] tvec = (trapToDebug ? {20'd0, debugTVec} : notDebugTVec);
	wire _io_eret_T = insn_call | insn_break;
	wire exception = _io_eret_T | io_exception;
	wire [1:0] _T_255 = insn_ret + insn_call;
	wire [1:0] _T_257 = insn_break + io_exception;
	wire [2:0] _T_259 = _T_255 + _T_257;
	wire _T_263 = ~reset;
	wire _GEN_46 = ((insn_wfi & _io_interrupt_T) & _io_decode_0_read_illegal_T_16) | reg_wfi;
	wire _GEN_48 = (io_retire | exception) | reg_singleStepped;
	wire [31:0] _epc_T = ~io_pc;
	wire [31:0] _epc_T_1 = _epc_T | 32'h00000001;
	wire [31:0] epc = ~_epc_T_1;
	wire [1:0] _reg_dcsr_cause_T = (causeIsDebugTrigger ? 2'h2 : 2'h1);
	wire [1:0] _reg_dcsr_cause_T_1 = (causeIsDebugInt ? 2'h3 : _reg_dcsr_cause_T);
	wire [2:0] _reg_dcsr_cause_T_2 = (reg_singleStepped ? 3'h4 : {1'd0, _reg_dcsr_cause_T_1});
	wire _GEN_51 = _io_decode_0_read_illegal_T_16 | reg_debug;
	wire [31:0] _GEN_52 = (_io_decode_0_read_illegal_T_16 ? epc : reg_dpc);
	wire [1:0] _GEN_73 = {1'd0, reg_mstatus_spp};
	wire _GEN_145 = (trapToDebug ? _GEN_51 : reg_debug);
	wire [31:0] _GEN_146 = (trapToDebug ? _GEN_52 : reg_dpc);
	wire [1:0] _GEN_170 = (trapToDebug ? {1'd0, reg_mstatus_spp} : _GEN_73);
	wire [31:0] _GEN_174 = (trapToDebug ? reg_mepc : epc);
	wire [31:0] _GEN_175 = (trapToDebug ? reg_mcause : cause);
	wire [31:0] _GEN_176 = (trapToDebug ? reg_mtval : io_tval);
	wire _GEN_178 = (trapToDebug ? reg_mstatus_mpie : reg_mstatus_mie);
	wire _GEN_180 = trapToDebug & reg_mstatus_mie;
	wire _GEN_182 = (exception ? _GEN_145 : reg_debug);
	wire [31:0] _GEN_183 = (exception ? _GEN_146 : reg_dpc);
	wire [1:0] _GEN_207 = (exception ? _GEN_170 : {1'd0, reg_mstatus_spp});
	wire [31:0] _GEN_211 = (exception ? _GEN_174 : reg_mepc);
	wire [31:0] _GEN_212 = (exception ? _GEN_175 : reg_mcause);
	wire [31:0] _GEN_213 = (exception ? _GEN_176 : reg_mtval);
	wire _GEN_215 = (exception ? _GEN_178 : reg_mstatus_mpie);
	wire _GEN_217 = (exception ? _GEN_180 : reg_mstatus_mie);
	wire [31:0] _GEN_239 = (io_rw_addr[10] & io_rw_addr[7] ? _T_28 : _T_22);
	wire _GEN_241 = (io_rw_addr[10] & io_rw_addr[7] ? _GEN_217 : reg_mstatus_mpie);
	wire _GEN_242 = (io_rw_addr[10] & io_rw_addr[7] ? _GEN_215 : 1'h1);
	wire _GEN_273 = (insn_ret ? _GEN_241 : _GEN_217);
	wire _GEN_274 = (insn_ret ? _GEN_242 : _GEN_215);
	reg io_status_cease_r;
	wire _GEN_279 = insn_cease | io_status_cease_r;
	wire [31:0] _io_rw_rdata_T_1 = (decoded_1 ? _T_16 : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_2 = (decoded_2 ? reg_bp_0_address : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_4 = (decoded_4 ? reg_misa : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_5 = (decoded_5 ? read_mstatus : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_6 = (decoded_6 ? read_mtvec : 32'h00000000);
	wire [15:0] _io_rw_rdata_T_7 = (decoded_7 ? read_mip : 16'h0000);
	wire [31:0] _io_rw_rdata_T_8 = (decoded_8 ? reg_mie : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_9 = (decoded_9 ? reg_mscratch : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_10 = (decoded_10 ? _T_22 : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_11 = (decoded_11 ? reg_mtval : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_12 = (decoded_12 ? reg_mcause : 32'h00000000);
	wire _io_rw_rdata_T_13 = decoded_13 & io_hartid;
	wire [31:0] _io_rw_rdata_T_14 = (decoded_14 ? _T_23 : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_15 = (decoded_15 ? _T_28 : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_16 = (decoded_16 ? reg_dscratch : 32'h00000000);
	wire [2:0] _io_rw_rdata_T_17 = (decoded_17 ? reg_mcountinhibit : 3'h0);
	wire [63:0] _io_rw_rdata_T_18 = (decoded_18 ? value_1 : 64'h0000000000000000);
	wire [63:0] _io_rw_rdata_T_19 = (decoded_19 ? value : 64'h0000000000000000);
	wire [31:0] _io_rw_rdata_T_107 = (decoded_107 ? value_1[63:32] : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_108 = (decoded_108 ? value[63:32] : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_109 = (decoded_109 ? _T_64 : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_110 = (decoded_110 ? _T_69 : 32'h00000000);
	wire [29:0] _io_rw_rdata_T_113 = (decoded_113 ? reg_pmp_0_addr : 30'h00000000);
	wire [29:0] _io_rw_rdata_T_114 = (decoded_114 ? reg_pmp_1_addr : 30'h00000000);
	wire [29:0] _io_rw_rdata_T_115 = (decoded_115 ? reg_pmp_2_addr : 30'h00000000);
	wire [29:0] _io_rw_rdata_T_116 = (decoded_116 ? reg_pmp_3_addr : 30'h00000000);
	wire [29:0] _io_rw_rdata_T_117 = (decoded_117 ? reg_pmp_4_addr : 30'h00000000);
	wire [29:0] _io_rw_rdata_T_118 = (decoded_118 ? reg_pmp_5_addr : 30'h00000000);
	wire [29:0] _io_rw_rdata_T_119 = (decoded_119 ? reg_pmp_6_addr : 30'h00000000);
	wire [29:0] _io_rw_rdata_T_120 = (decoded_120 ? reg_pmp_7_addr : 30'h00000000);
	wire [31:0] _io_rw_rdata_T_129 = (decoded_129 ? reg_custom_0 : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_130 = (decoded_130 ? 32'h00000001 : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_132 = (decoded_132 ? 32'h20181004 : 32'h00000000);
	wire [31:0] _io_rw_rdata_T_134 = _io_rw_rdata_T_1 | _io_rw_rdata_T_2;
	wire [31:0] _io_rw_rdata_T_136 = _io_rw_rdata_T_134 | _io_rw_rdata_T_4;
	wire [31:0] _io_rw_rdata_T_137 = _io_rw_rdata_T_136 | _io_rw_rdata_T_5;
	wire [31:0] _io_rw_rdata_T_138 = _io_rw_rdata_T_137 | _io_rw_rdata_T_6;
	wire [31:0] _GEN_592 = {16'd0, _io_rw_rdata_T_7};
	wire [31:0] _io_rw_rdata_T_139 = _io_rw_rdata_T_138 | _GEN_592;
	wire [31:0] _io_rw_rdata_T_140 = _io_rw_rdata_T_139 | _io_rw_rdata_T_8;
	wire [31:0] _io_rw_rdata_T_141 = _io_rw_rdata_T_140 | _io_rw_rdata_T_9;
	wire [31:0] _io_rw_rdata_T_142 = _io_rw_rdata_T_141 | _io_rw_rdata_T_10;
	wire [31:0] _io_rw_rdata_T_143 = _io_rw_rdata_T_142 | _io_rw_rdata_T_11;
	wire [31:0] _io_rw_rdata_T_144 = _io_rw_rdata_T_143 | _io_rw_rdata_T_12;
	wire [31:0] _GEN_593 = {31'd0, _io_rw_rdata_T_13};
	wire [31:0] _io_rw_rdata_T_145 = _io_rw_rdata_T_144 | _GEN_593;
	wire [31:0] _io_rw_rdata_T_146 = _io_rw_rdata_T_145 | _io_rw_rdata_T_14;
	wire [31:0] _io_rw_rdata_T_147 = _io_rw_rdata_T_146 | _io_rw_rdata_T_15;
	wire [31:0] _io_rw_rdata_T_148 = _io_rw_rdata_T_147 | _io_rw_rdata_T_16;
	wire [31:0] _GEN_594 = {29'd0, _io_rw_rdata_T_17};
	wire [31:0] _io_rw_rdata_T_149 = _io_rw_rdata_T_148 | _GEN_594;
	wire [63:0] _GEN_595 = {32'd0, _io_rw_rdata_T_149};
	wire [63:0] _io_rw_rdata_T_150 = _GEN_595 | _io_rw_rdata_T_18;
	wire [63:0] _io_rw_rdata_T_151 = _io_rw_rdata_T_150 | _io_rw_rdata_T_19;
	wire [63:0] _GEN_596 = {32'd0, _io_rw_rdata_T_107};
	wire [63:0] _io_rw_rdata_T_239 = _io_rw_rdata_T_151 | _GEN_596;
	wire [63:0] _GEN_597 = {32'd0, _io_rw_rdata_T_108};
	wire [63:0] _io_rw_rdata_T_240 = _io_rw_rdata_T_239 | _GEN_597;
	wire [63:0] _GEN_598 = {32'd0, _io_rw_rdata_T_109};
	wire [63:0] _io_rw_rdata_T_241 = _io_rw_rdata_T_240 | _GEN_598;
	wire [63:0] _GEN_599 = {32'd0, _io_rw_rdata_T_110};
	wire [63:0] _io_rw_rdata_T_242 = _io_rw_rdata_T_241 | _GEN_599;
	wire [63:0] _GEN_600 = {34'd0, _io_rw_rdata_T_113};
	wire [63:0] _io_rw_rdata_T_245 = _io_rw_rdata_T_242 | _GEN_600;
	wire [63:0] _GEN_601 = {34'd0, _io_rw_rdata_T_114};
	wire [63:0] _io_rw_rdata_T_246 = _io_rw_rdata_T_245 | _GEN_601;
	wire [63:0] _GEN_602 = {34'd0, _io_rw_rdata_T_115};
	wire [63:0] _io_rw_rdata_T_247 = _io_rw_rdata_T_246 | _GEN_602;
	wire [63:0] _GEN_603 = {34'd0, _io_rw_rdata_T_116};
	wire [63:0] _io_rw_rdata_T_248 = _io_rw_rdata_T_247 | _GEN_603;
	wire [63:0] _GEN_604 = {34'd0, _io_rw_rdata_T_117};
	wire [63:0] _io_rw_rdata_T_249 = _io_rw_rdata_T_248 | _GEN_604;
	wire [63:0] _GEN_605 = {34'd0, _io_rw_rdata_T_118};
	wire [63:0] _io_rw_rdata_T_250 = _io_rw_rdata_T_249 | _GEN_605;
	wire [63:0] _GEN_606 = {34'd0, _io_rw_rdata_T_119};
	wire [63:0] _io_rw_rdata_T_251 = _io_rw_rdata_T_250 | _GEN_606;
	wire [63:0] _GEN_607 = {34'd0, _io_rw_rdata_T_120};
	wire [63:0] _io_rw_rdata_T_252 = _io_rw_rdata_T_251 | _GEN_607;
	wire [63:0] _GEN_608 = {32'd0, _io_rw_rdata_T_129};
	wire [63:0] _io_rw_rdata_T_261 = _io_rw_rdata_T_252 | _GEN_608;
	wire [63:0] _GEN_609 = {32'd0, _io_rw_rdata_T_130};
	wire [63:0] _io_rw_rdata_T_262 = _io_rw_rdata_T_261 | _GEN_609;
	wire [63:0] _GEN_610 = {32'd0, _io_rw_rdata_T_132};
	wire [63:0] _io_rw_rdata_T_264 = _io_rw_rdata_T_262 | _GEN_610;
	wire _T_407 = io_rw_cmd == 3'h5;
	wire _T_408 = io_rw_cmd == 3'h6;
	wire _T_409 = io_rw_cmd == 3'h7;
	wire csr_wen = (_T_408 | _T_409) | _T_407;
	wire [104:0] _new_mstatus_WIRE = {73'd0, wdata};
	wire new_mstatus_mie = _new_mstatus_WIRE[3];
	wire new_mstatus_mpie = _new_mstatus_WIRE[7];
	wire f = wdata[5];
	wire [31:0] _reg_misa_T = ~wdata;
	wire _reg_misa_T_1 = ~f;
	wire [3:0] _reg_misa_T_2 = {_reg_misa_T_1, 3'h0};
	wire [31:0] _GEN_611 = {28'd0, _reg_misa_T_2};
	wire [31:0] _reg_misa_T_3 = _reg_misa_T | _GEN_611;
	wire [31:0] _reg_misa_T_4 = ~_reg_misa_T_3;
	wire [31:0] _reg_misa_T_5 = _reg_misa_T_4 & 32'h00001005;
	wire [31:0] _reg_misa_T_7 = reg_misa & 32'hffffeffa;
	wire [31:0] _reg_misa_T_8 = _reg_misa_T_5 | _reg_misa_T_7;
	wire [31:0] _reg_mie_T = wdata & 32'h00000888;
	wire [31:0] _reg_mepc_T_1 = _reg_misa_T | 32'h00000001;
	wire [31:0] _reg_mepc_T_2 = ~_reg_mepc_T_1;
	wire [31:0] _reg_mcause_T = wdata & 32'h8000000f;
	wire [31:0] _reg_mcountinhibit_T_1 = wdata & 32'hfffffffd;
	wire [31:0] _GEN_295 = (decoded_17 ? _reg_mcountinhibit_T_1 : {29'd0, reg_mcountinhibit});
	wire [63:0] _T_2007 = {value_1[63:32], wdata};
	wire [63:0] _GEN_296 = (decoded_18 ? _T_2007 : {57'd0, _GEN_2});
	wire [63:0] _T_2010 = {wdata, value_1[31:0]};
	wire [63:0] _GEN_298 = (decoded_107 ? _T_2010 : _GEN_296);
	wire [63:0] _T_2012 = {value[63:32], wdata};
	wire [63:0] _GEN_300 = (decoded_19 ? _T_2012 : {57'd0, _GEN_0});
	wire [63:0] _T_2015 = {wdata, value[31:0]};
	wire [63:0] _GEN_302 = (decoded_108 ? _T_2015 : _GEN_300);
	wire new_dcsr_ebreakm = wdata[15];
	wire [31:0] _newBPC_T_2 = (io_rw_cmd[1] ? _T_16 : 32'h00000000);
	wire [31:0] _newBPC_T_3 = _newBPC_T_2 | io_rw_wdata;
	wire [31:0] _newBPC_T_8 = _newBPC_T_3 & _wdata_T_6;
	wire newBPC_action = _newBPC_T_8[12];
	wire newBPC_dmode = _newBPC_T_8[27];
	wire dMode = newBPC_dmode & reg_debug;
	wire _GEN_310 = dMode & newBPC_action;
	wire newCfg_r = wdata[0];
	wire newCfg_w = wdata[1];
	wire newCfg_x = wdata[2];
	wire [1:0] newCfg_a = wdata[4:3];
	wire newCfg_l = wdata[7];
	wire _T_2033 = ~reg_pmp_1_cfg_a[1] & reg_pmp_1_cfg_a[0];
	wire _T_2035 = reg_pmp_0_cfg_l | (reg_pmp_1_cfg_l & _T_2033);
	wire [31:0] _GEN_381 = (decoded_113 & ~_T_2035 ? wdata : {2'd0, reg_pmp_0_addr});
	wire newCfg_1_r = wdata[8];
	wire newCfg_1_w = wdata[9];
	wire newCfg_1_x = wdata[10];
	wire [1:0] newCfg_1_a = wdata[12:11];
	wire newCfg_1_l = wdata[15];
	wire _T_2043 = ~reg_pmp_2_cfg_a[1] & reg_pmp_2_cfg_a[0];
	wire _T_2045 = reg_pmp_1_cfg_l | (reg_pmp_2_cfg_l & _T_2043);
	wire [31:0] _GEN_388 = (decoded_114 & ~_T_2045 ? wdata : {2'd0, reg_pmp_1_addr});
	wire newCfg_2_r = wdata[16];
	wire newCfg_2_w = wdata[17];
	wire newCfg_2_x = wdata[18];
	wire [1:0] newCfg_2_a = wdata[20:19];
	wire newCfg_2_l = wdata[23];
	wire _T_2053 = ~reg_pmp_3_cfg_a[1] & reg_pmp_3_cfg_a[0];
	wire _T_2055 = reg_pmp_2_cfg_l | (reg_pmp_3_cfg_l & _T_2053);
	wire [31:0] _GEN_395 = (decoded_115 & ~_T_2055 ? wdata : {2'd0, reg_pmp_2_addr});
	wire newCfg_3_r = wdata[24];
	wire newCfg_3_w = wdata[25];
	wire newCfg_3_x = wdata[26];
	wire [1:0] newCfg_3_a = wdata[28:27];
	wire newCfg_3_l = wdata[31];
	wire _T_2063 = ~reg_pmp_4_cfg_a[1] & reg_pmp_4_cfg_a[0];
	wire _T_2065 = reg_pmp_3_cfg_l | (reg_pmp_4_cfg_l & _T_2063);
	wire [31:0] _GEN_402 = (decoded_116 & ~_T_2065 ? wdata : {2'd0, reg_pmp_3_addr});
	wire _T_2073 = ~reg_pmp_5_cfg_a[1] & reg_pmp_5_cfg_a[0];
	wire _T_2075 = reg_pmp_4_cfg_l | (reg_pmp_5_cfg_l & _T_2073);
	wire [31:0] _GEN_409 = (decoded_117 & ~_T_2075 ? wdata : {2'd0, reg_pmp_4_addr});
	wire _T_2083 = ~reg_pmp_6_cfg_a[1] & reg_pmp_6_cfg_a[0];
	wire _T_2085 = reg_pmp_5_cfg_l | (reg_pmp_6_cfg_l & _T_2083);
	wire [31:0] _GEN_416 = (decoded_118 & ~_T_2085 ? wdata : {2'd0, reg_pmp_5_addr});
	wire _T_2093 = ~reg_pmp_7_cfg_a[1] & reg_pmp_7_cfg_a[0];
	wire _T_2095 = reg_pmp_6_cfg_l | (reg_pmp_7_cfg_l & _T_2093);
	wire [31:0] _GEN_423 = (decoded_119 & ~_T_2095 ? wdata : {2'd0, reg_pmp_6_addr});
	wire _T_2105 = reg_pmp_7_cfg_l | (reg_pmp_7_cfg_l & _T_2093);
	wire [31:0] _GEN_430 = (decoded_120 & ~_T_2105 ? wdata : {2'd0, reg_pmp_7_addr});
	wire [31:0] _reg_custom_0_T = wdata & 32'h00000008;
	wire [31:0] _reg_custom_0_T_2 = reg_custom_0 & 32'hfffffff7;
	wire [31:0] _reg_custom_0_T_3 = _reg_custom_0_T | _reg_custom_0_T_2;
	wire [31:0] _GEN_449 = (csr_wen ? _GEN_295 : {29'd0, reg_mcountinhibit});
	wire [63:0] _GEN_450 = (csr_wen ? _GEN_298 : {57'd0, _GEN_2});
	wire [63:0] _GEN_452 = (csr_wen ? _GEN_302 : {57'd0, _GEN_0});
	wire [31:0] _GEN_497 = (csr_wen ? _GEN_381 : {2'd0, reg_pmp_0_addr});
	wire [31:0] _GEN_504 = (csr_wen ? _GEN_388 : {2'd0, reg_pmp_1_addr});
	wire [31:0] _GEN_511 = (csr_wen ? _GEN_395 : {2'd0, reg_pmp_2_addr});
	wire [31:0] _GEN_518 = (csr_wen ? _GEN_402 : {2'd0, reg_pmp_3_addr});
	wire [31:0] _GEN_525 = (csr_wen ? _GEN_409 : {2'd0, reg_pmp_4_addr});
	wire [31:0] _GEN_532 = (csr_wen ? _GEN_416 : {2'd0, reg_pmp_5_addr});
	wire [31:0] _GEN_539 = (csr_wen ? _GEN_423 : {2'd0, reg_pmp_6_addr});
	wire [31:0] _GEN_546 = (csr_wen ? _GEN_430 : {2'd0, reg_pmp_7_addr});
	assign io_rw_rdata = _io_rw_rdata_T_264[31:0];
	assign io_decode_0_fp_illegal = (io_status_fs == 2'h0) | ~reg_misa[5];
	assign io_decode_0_fp_csr = 1'h0;
	assign io_decode_0_read_illegal = _io_decode_0_read_illegal_T_18 | _io_decode_0_read_illegal_T_21;
	assign io_decode_0_write_illegal = &addr_1[11:10];
	assign io_decode_0_write_flush = ~((io_decode_0_write_flush_addr_m >= 12'h340) & (io_decode_0_write_flush_addr_m <= 12'h343));
	assign io_decode_0_system_illegal = ((is_ret & addr_1[10]) & addr_1[7]) & _io_decode_0_read_illegal_T_16;
	assign io_csr_stall = reg_wfi | io_status_cease;
	assign io_eret = (insn_call | insn_break) | insn_ret;
	assign io_singleStep = reg_dcsr_step & _io_decode_0_read_illegal_T_16;
	assign io_status_debug = reg_debug;
	assign io_status_cease = io_status_cease_r;
	assign io_status_wfi = reg_wfi;
	assign io_status_isa = reg_misa;
	assign io_status_dprv = 2'h3;
	assign io_status_dv = 1'h0;
	assign io_status_prv = 2'h3;
	assign io_status_v = 1'h0;
	assign io_status_sd = (&io_status_fs | &io_status_xs) | &io_status_vs;
	assign io_status_zero2 = 23'h000000;
	assign io_status_mpv = 1'h0;
	assign io_status_gva = reg_mstatus_gva;
	assign io_status_mbe = 1'h0;
	assign io_status_sbe = 1'h0;
	assign io_status_sxl = 2'h0;
	assign io_status_uxl = 2'h0;
	assign io_status_sd_rv32 = io_status_sd;
	assign io_status_zero1 = 8'h00;
	assign io_status_tsr = 1'h0;
	assign io_status_tw = 1'h0;
	assign io_status_tvm = 1'h0;
	assign io_status_mxr = 1'h0;
	assign io_status_sum = 1'h0;
	assign io_status_mprv = 1'h0;
	assign io_status_xs = 2'h0;
	assign io_status_fs = 2'h0;
	assign io_status_mpp = 2'h3;
	assign io_status_vs = 2'h0;
	assign io_status_spp = reg_mstatus_spp;
	assign io_status_mpie = reg_mstatus_mpie;
	assign io_status_ube = 1'h0;
	assign io_status_spie = 1'h0;
	assign io_status_upie = 1'h0;
	assign io_status_mie = reg_mstatus_mie;
	assign io_status_hie = 1'h0;
	assign io_status_sie = 1'h0;
	assign io_status_uie = 1'h0;
	assign io_evec = (insn_ret ? _GEN_239 : tvec);
	assign io_time = value_1[31:0];
	assign io_interrupt = ((anyInterrupt & ~io_singleStep) | reg_singleStepped) & ~(reg_debug | io_status_cease);
	assign io_interrupt_cause = 32'h80000000 + _GEN_41;
	assign io_bp_0_control_action = reg_bp_0_control_action;
	assign io_bp_0_control_tmatch = reg_bp_0_control_tmatch;
	assign io_bp_0_control_x = reg_bp_0_control_x;
	assign io_bp_0_control_w = reg_bp_0_control_w;
	assign io_bp_0_control_r = reg_bp_0_control_r;
	assign io_bp_0_address = reg_bp_0_address;
	assign io_pmp_0_cfg_l = reg_pmp_0_cfg_l;
	assign io_pmp_0_cfg_a = reg_pmp_0_cfg_a;
	assign io_pmp_0_cfg_x = reg_pmp_0_cfg_x;
	assign io_pmp_0_cfg_w = reg_pmp_0_cfg_w;
	assign io_pmp_0_cfg_r = reg_pmp_0_cfg_r;
	assign io_pmp_0_addr = reg_pmp_0_addr;
	assign io_pmp_0_mask = _pmp_mask_T_4[31:0];
	assign io_pmp_1_cfg_l = reg_pmp_1_cfg_l;
	assign io_pmp_1_cfg_a = reg_pmp_1_cfg_a;
	assign io_pmp_1_cfg_x = reg_pmp_1_cfg_x;
	assign io_pmp_1_cfg_w = reg_pmp_1_cfg_w;
	assign io_pmp_1_cfg_r = reg_pmp_1_cfg_r;
	assign io_pmp_1_addr = reg_pmp_1_addr;
	assign io_pmp_1_mask = _pmp_mask_T_9[31:0];
	assign io_pmp_2_cfg_l = reg_pmp_2_cfg_l;
	assign io_pmp_2_cfg_a = reg_pmp_2_cfg_a;
	assign io_pmp_2_cfg_x = reg_pmp_2_cfg_x;
	assign io_pmp_2_cfg_w = reg_pmp_2_cfg_w;
	assign io_pmp_2_cfg_r = reg_pmp_2_cfg_r;
	assign io_pmp_2_addr = reg_pmp_2_addr;
	assign io_pmp_2_mask = _pmp_mask_T_14[31:0];
	assign io_pmp_3_cfg_l = reg_pmp_3_cfg_l;
	assign io_pmp_3_cfg_a = reg_pmp_3_cfg_a;
	assign io_pmp_3_cfg_x = reg_pmp_3_cfg_x;
	assign io_pmp_3_cfg_w = reg_pmp_3_cfg_w;
	assign io_pmp_3_cfg_r = reg_pmp_3_cfg_r;
	assign io_pmp_3_addr = reg_pmp_3_addr;
	assign io_pmp_3_mask = _pmp_mask_T_19[31:0];
	assign io_pmp_4_cfg_l = reg_pmp_4_cfg_l;
	assign io_pmp_4_cfg_a = reg_pmp_4_cfg_a;
	assign io_pmp_4_cfg_x = reg_pmp_4_cfg_x;
	assign io_pmp_4_cfg_w = reg_pmp_4_cfg_w;
	assign io_pmp_4_cfg_r = reg_pmp_4_cfg_r;
	assign io_pmp_4_addr = reg_pmp_4_addr;
	assign io_pmp_4_mask = _pmp_mask_T_24[31:0];
	assign io_pmp_5_cfg_l = reg_pmp_5_cfg_l;
	assign io_pmp_5_cfg_a = reg_pmp_5_cfg_a;
	assign io_pmp_5_cfg_x = reg_pmp_5_cfg_x;
	assign io_pmp_5_cfg_w = reg_pmp_5_cfg_w;
	assign io_pmp_5_cfg_r = reg_pmp_5_cfg_r;
	assign io_pmp_5_addr = reg_pmp_5_addr;
	assign io_pmp_5_mask = _pmp_mask_T_29[31:0];
	assign io_pmp_6_cfg_l = reg_pmp_6_cfg_l;
	assign io_pmp_6_cfg_a = reg_pmp_6_cfg_a;
	assign io_pmp_6_cfg_x = reg_pmp_6_cfg_x;
	assign io_pmp_6_cfg_w = reg_pmp_6_cfg_w;
	assign io_pmp_6_cfg_r = reg_pmp_6_cfg_r;
	assign io_pmp_6_addr = reg_pmp_6_addr;
	assign io_pmp_6_mask = _pmp_mask_T_34[31:0];
	assign io_pmp_7_cfg_l = reg_pmp_7_cfg_l;
	assign io_pmp_7_cfg_a = reg_pmp_7_cfg_a;
	assign io_pmp_7_cfg_x = reg_pmp_7_cfg_x;
	assign io_pmp_7_cfg_w = reg_pmp_7_cfg_w;
	assign io_pmp_7_cfg_r = reg_pmp_7_cfg_r;
	assign io_pmp_7_addr = reg_pmp_7_addr;
	assign io_pmp_7_mask = _pmp_mask_T_39[31:0];
	assign io_inhibit_cycle = reg_mcountinhibit[0];
	assign io_trace_0_valid = (io_retire > 1'h0) | io_trace_0_exception;
	assign io_trace_0_iaddr = io_pc;
	assign io_trace_0_insn = io_inst_0;
	assign io_trace_0_exception = _io_eret_T | io_exception;
	assign io_customCSRs_0_value = reg_custom_0;
	always @(posedge clock) begin
		if (reset)
			reg_mstatus_gva <= 1'h0;
		else if (exception)
			if (!trapToDebug)
				reg_mstatus_gva <= io_gva;
		if (reset)
			reg_mstatus_spp <= 1'h0;
		else
			reg_mstatus_spp <= _GEN_207[0];
		if (reset)
			reg_mstatus_mpie <= 1'h0;
		else if (csr_wen) begin
			if (decoded_5)
				reg_mstatus_mpie <= new_mstatus_mpie;
			else
				reg_mstatus_mpie <= _GEN_274;
		end
		else
			reg_mstatus_mpie <= _GEN_274;
		if (reset)
			reg_mstatus_mie <= 1'h0;
		else if (csr_wen) begin
			if (decoded_5)
				reg_mstatus_mie <= new_mstatus_mie;
			else
				reg_mstatus_mie <= _GEN_273;
		end
		else
			reg_mstatus_mie <= _GEN_273;
		if (reset)
			reg_dcsr_ebreakm <= 1'h0;
		else if (csr_wen)
			if (decoded_14)
				reg_dcsr_ebreakm <= new_dcsr_ebreakm;
		if (reset)
			reg_dcsr_cause <= 3'h0;
		else if (exception)
			if (trapToDebug)
				if (_io_decode_0_read_illegal_T_16)
					reg_dcsr_cause <= _reg_dcsr_cause_T_2;
		if (reset)
			reg_dcsr_step <= 1'h0;
		else if (csr_wen)
			if (decoded_14)
				reg_dcsr_step <= wdata[2];
		if (reset)
			reg_debug <= 1'h0;
		else if (insn_ret) begin
			if (io_rw_addr[10] & io_rw_addr[7])
				reg_debug <= 1'h0;
			else
				reg_debug <= _GEN_182;
		end
		else
			reg_debug <= _GEN_182;
		if (csr_wen) begin
			if (decoded_15)
				reg_dpc <= _reg_mepc_T_2;
			else
				reg_dpc <= _GEN_183;
		end
		else
			reg_dpc <= _GEN_183;
		if (csr_wen)
			if (decoded_16)
				reg_dscratch <= wdata;
		if (_io_interrupt_T)
			reg_singleStepped <= 1'h0;
		else
			reg_singleStepped <= _GEN_48;
		if (reset)
			reg_bp_0_control_dmode <= 1'h0;
		else if (csr_wen)
			if (~reg_bp_0_control_dmode | reg_debug)
				if (decoded_1)
					reg_bp_0_control_dmode <= dMode;
		if (reset)
			reg_bp_0_control_action <= 1'h0;
		else if (csr_wen)
			if (~reg_bp_0_control_dmode | reg_debug)
				if (decoded_1)
					reg_bp_0_control_action <= _GEN_310;
		if (csr_wen)
			if (~reg_bp_0_control_dmode | reg_debug)
				if (decoded_1)
					reg_bp_0_control_tmatch <= wdata[8:7];
		if (reset)
			reg_bp_0_control_x <= 1'h0;
		else if (csr_wen)
			if (~reg_bp_0_control_dmode | reg_debug)
				if (decoded_1)
					reg_bp_0_control_x <= wdata[2];
		if (reset)
			reg_bp_0_control_w <= 1'h0;
		else if (csr_wen)
			if (~reg_bp_0_control_dmode | reg_debug)
				if (decoded_1)
					reg_bp_0_control_w <= wdata[1];
		if (reset)
			reg_bp_0_control_r <= 1'h0;
		else if (csr_wen)
			if (~reg_bp_0_control_dmode | reg_debug)
				if (decoded_1)
					reg_bp_0_control_r <= wdata[0];
		if (csr_wen)
			if (~reg_bp_0_control_dmode | reg_debug)
				if (decoded_2)
					reg_bp_0_address <= wdata;
		if (reset)
			reg_pmp_0_cfg_l <= 1'h0;
		else if (csr_wen)
			if (decoded_109 & ~reg_pmp_0_cfg_l)
				reg_pmp_0_cfg_l <= newCfg_l;
		if (reset)
			reg_pmp_0_cfg_a <= 2'h0;
		else if (csr_wen)
			if (decoded_109 & ~reg_pmp_0_cfg_l)
				reg_pmp_0_cfg_a <= newCfg_a;
		if (csr_wen)
			if (decoded_109 & ~reg_pmp_0_cfg_l)
				reg_pmp_0_cfg_x <= newCfg_x;
		if (csr_wen)
			if (decoded_109 & ~reg_pmp_0_cfg_l)
				reg_pmp_0_cfg_w <= newCfg_w & newCfg_r;
		if (csr_wen)
			if (decoded_109 & ~reg_pmp_0_cfg_l)
				reg_pmp_0_cfg_r <= newCfg_r;
		reg_pmp_0_addr <= _GEN_497[29:0];
		if (reset)
			reg_pmp_1_cfg_l <= 1'h0;
		else if (csr_wen)
			if (decoded_109 & ~reg_pmp_1_cfg_l)
				reg_pmp_1_cfg_l <= newCfg_1_l;
		if (reset)
			reg_pmp_1_cfg_a <= 2'h0;
		else if (csr_wen)
			if (decoded_109 & ~reg_pmp_1_cfg_l)
				reg_pmp_1_cfg_a <= newCfg_1_a;
		if (csr_wen)
			if (decoded_109 & ~reg_pmp_1_cfg_l)
				reg_pmp_1_cfg_x <= newCfg_1_x;
		if (csr_wen)
			if (decoded_109 & ~reg_pmp_1_cfg_l)
				reg_pmp_1_cfg_w <= newCfg_1_w & newCfg_1_r;
		if (csr_wen)
			if (decoded_109 & ~reg_pmp_1_cfg_l)
				reg_pmp_1_cfg_r <= newCfg_1_r;
		reg_pmp_1_addr <= _GEN_504[29:0];
		if (reset)
			reg_pmp_2_cfg_l <= 1'h0;
		else if (csr_wen)
			if (decoded_109 & ~reg_pmp_2_cfg_l)
				reg_pmp_2_cfg_l <= newCfg_2_l;
		if (reset)
			reg_pmp_2_cfg_a <= 2'h0;
		else if (csr_wen)
			if (decoded_109 & ~reg_pmp_2_cfg_l)
				reg_pmp_2_cfg_a <= newCfg_2_a;
		if (csr_wen)
			if (decoded_109 & ~reg_pmp_2_cfg_l)
				reg_pmp_2_cfg_x <= newCfg_2_x;
		if (csr_wen)
			if (decoded_109 & ~reg_pmp_2_cfg_l)
				reg_pmp_2_cfg_w <= newCfg_2_w & newCfg_2_r;
		if (csr_wen)
			if (decoded_109 & ~reg_pmp_2_cfg_l)
				reg_pmp_2_cfg_r <= newCfg_2_r;
		reg_pmp_2_addr <= _GEN_511[29:0];
		if (reset)
			reg_pmp_3_cfg_l <= 1'h0;
		else if (csr_wen)
			if (decoded_109 & ~reg_pmp_3_cfg_l)
				reg_pmp_3_cfg_l <= newCfg_3_l;
		if (reset)
			reg_pmp_3_cfg_a <= 2'h0;
		else if (csr_wen)
			if (decoded_109 & ~reg_pmp_3_cfg_l)
				reg_pmp_3_cfg_a <= newCfg_3_a;
		if (csr_wen)
			if (decoded_109 & ~reg_pmp_3_cfg_l)
				reg_pmp_3_cfg_x <= newCfg_3_x;
		if (csr_wen)
			if (decoded_109 & ~reg_pmp_3_cfg_l)
				reg_pmp_3_cfg_w <= newCfg_3_w & newCfg_3_r;
		if (csr_wen)
			if (decoded_109 & ~reg_pmp_3_cfg_l)
				reg_pmp_3_cfg_r <= newCfg_3_r;
		reg_pmp_3_addr <= _GEN_518[29:0];
		if (reset)
			reg_pmp_4_cfg_l <= 1'h0;
		else if (csr_wen)
			if (decoded_110 & ~reg_pmp_4_cfg_l)
				reg_pmp_4_cfg_l <= newCfg_l;
		if (reset)
			reg_pmp_4_cfg_a <= 2'h0;
		else if (csr_wen)
			if (decoded_110 & ~reg_pmp_4_cfg_l)
				reg_pmp_4_cfg_a <= newCfg_a;
		if (csr_wen)
			if (decoded_110 & ~reg_pmp_4_cfg_l)
				reg_pmp_4_cfg_x <= newCfg_x;
		if (csr_wen)
			if (decoded_110 & ~reg_pmp_4_cfg_l)
				reg_pmp_4_cfg_w <= newCfg_w & newCfg_r;
		if (csr_wen)
			if (decoded_110 & ~reg_pmp_4_cfg_l)
				reg_pmp_4_cfg_r <= newCfg_r;
		reg_pmp_4_addr <= _GEN_525[29:0];
		if (reset)
			reg_pmp_5_cfg_l <= 1'h0;
		else if (csr_wen)
			if (decoded_110 & ~reg_pmp_5_cfg_l)
				reg_pmp_5_cfg_l <= newCfg_1_l;
		if (reset)
			reg_pmp_5_cfg_a <= 2'h0;
		else if (csr_wen)
			if (decoded_110 & ~reg_pmp_5_cfg_l)
				reg_pmp_5_cfg_a <= newCfg_1_a;
		if (csr_wen)
			if (decoded_110 & ~reg_pmp_5_cfg_l)
				reg_pmp_5_cfg_x <= newCfg_1_x;
		if (csr_wen)
			if (decoded_110 & ~reg_pmp_5_cfg_l)
				reg_pmp_5_cfg_w <= newCfg_1_w & newCfg_1_r;
		if (csr_wen)
			if (decoded_110 & ~reg_pmp_5_cfg_l)
				reg_pmp_5_cfg_r <= newCfg_1_r;
		reg_pmp_5_addr <= _GEN_532[29:0];
		if (reset)
			reg_pmp_6_cfg_l <= 1'h0;
		else if (csr_wen)
			if (decoded_110 & ~reg_pmp_6_cfg_l)
				reg_pmp_6_cfg_l <= newCfg_2_l;
		if (reset)
			reg_pmp_6_cfg_a <= 2'h0;
		else if (csr_wen)
			if (decoded_110 & ~reg_pmp_6_cfg_l)
				reg_pmp_6_cfg_a <= newCfg_2_a;
		if (csr_wen)
			if (decoded_110 & ~reg_pmp_6_cfg_l)
				reg_pmp_6_cfg_x <= newCfg_2_x;
		if (csr_wen)
			if (decoded_110 & ~reg_pmp_6_cfg_l)
				reg_pmp_6_cfg_w <= newCfg_2_w & newCfg_2_r;
		if (csr_wen)
			if (decoded_110 & ~reg_pmp_6_cfg_l)
				reg_pmp_6_cfg_r <= newCfg_2_r;
		reg_pmp_6_addr <= _GEN_539[29:0];
		if (reset)
			reg_pmp_7_cfg_l <= 1'h0;
		else if (csr_wen)
			if (decoded_110 & ~reg_pmp_7_cfg_l)
				reg_pmp_7_cfg_l <= newCfg_3_l;
		if (reset)
			reg_pmp_7_cfg_a <= 2'h0;
		else if (csr_wen)
			if (decoded_110 & ~reg_pmp_7_cfg_l)
				reg_pmp_7_cfg_a <= newCfg_3_a;
		if (csr_wen)
			if (decoded_110 & ~reg_pmp_7_cfg_l)
				reg_pmp_7_cfg_x <= newCfg_3_x;
		if (csr_wen)
			if (decoded_110 & ~reg_pmp_7_cfg_l)
				reg_pmp_7_cfg_w <= newCfg_3_w & newCfg_3_r;
		if (csr_wen)
			if (decoded_110 & ~reg_pmp_7_cfg_l)
				reg_pmp_7_cfg_r <= newCfg_3_r;
		reg_pmp_7_addr <= _GEN_546[29:0];
		if (csr_wen)
			if (decoded_8)
				reg_mie <= _reg_mie_T;
		if (csr_wen) begin
			if (decoded_10)
				reg_mepc <= _reg_mepc_T_2;
			else
				reg_mepc <= _GEN_211;
		end
		else
			reg_mepc <= _GEN_211;
		if (reset)
			reg_mcause <= 32'h00000000;
		else if (csr_wen) begin
			if (decoded_12)
				reg_mcause <= _reg_mcause_T;
			else
				reg_mcause <= _GEN_212;
		end
		else
			reg_mcause <= _GEN_212;
		if (csr_wen) begin
			if (decoded_11)
				reg_mtval <= wdata;
			else
				reg_mtval <= _GEN_213;
		end
		else
			reg_mtval <= _GEN_213;
		if (csr_wen)
			if (decoded_9)
				reg_mscratch <= wdata;
		if (reset)
			reg_mtvec <= 32'h00000000;
		else if (csr_wen)
			if (decoded_6)
				reg_mtvec <= wdata;
		if (reset)
			reg_mcountinhibit <= 3'h0;
		else
			reg_mcountinhibit <= _GEN_449[2:0];
		if (reset)
			small_ <= 6'h00;
		else
			small_ <= _GEN_452[5:0];
		if (reset)
			large_ <= 58'h000000000000000;
		else if (csr_wen) begin
			if (decoded_108)
				large_ <= _T_2015[63:6];
			else if (decoded_19)
				large_ <= _T_2012[63:6];
			else
				large_ <= _GEN_1;
		end
		else
			large_ <= _GEN_1;
		if (reset)
			reg_misa <= 32'h40801105;
		else if (csr_wen)
			if (decoded_4)
				if (~io_pc[1] | wdata[2])
					reg_misa <= _reg_misa_T_8;
		if (reset)
			reg_custom_0 <= 32'h00000008;
		else if (csr_wen)
			if (decoded_129)
				reg_custom_0 <= _reg_custom_0_T_3;
		if (reset)
			io_status_cease_r <= 1'h0;
		else
			io_status_cease_r <= _GEN_279;
	end
	always @(posedge io_ungated_clock) begin
		if (reset)
			reg_wfi <= 1'h0;
		else if ((|pending_interrupts | io_interrupts_debug) | exception)
			reg_wfi <= 1'h0;
		else
			reg_wfi <= _GEN_46;
		if (reset)
			small_1 <= 6'h00;
		else
			small_1 <= _GEN_450[5:0];
		if (reset)
			large_1 <= 58'h000000000000000;
		else if (csr_wen) begin
			if (decoded_107)
				large_1 <= _T_2010[63:6];
			else if (decoded_18)
				large_1 <= _T_2007[63:6];
			else
				large_1 <= _GEN_3;
		end
		else
			large_1 <= _GEN_3;
	end
endmodule
module BreakpointUnit (
	io_status_debug,
	io_bp_0_control_action,
	io_bp_0_control_tmatch,
	io_bp_0_control_x,
	io_bp_0_control_w,
	io_bp_0_control_r,
	io_bp_0_address,
	io_pc,
	io_ea,
	io_xcpt_if,
	io_xcpt_ld,
	io_xcpt_st,
	io_debug_if,
	io_debug_ld,
	io_debug_st
);
	input io_status_debug;
	input io_bp_0_control_action;
	input [1:0] io_bp_0_control_tmatch;
	input io_bp_0_control_x;
	input io_bp_0_control_w;
	input io_bp_0_control_r;
	input [31:0] io_bp_0_address;
	input [31:0] io_pc;
	input [31:0] io_ea;
	output wire io_xcpt_if;
	output wire io_xcpt_ld;
	output wire io_xcpt_st;
	output wire io_debug_if;
	output wire io_debug_ld;
	output wire io_debug_st;
	wire en = ~io_status_debug;
	wire _r_T_4 = (io_ea >= io_bp_0_address) ^ io_bp_0_control_tmatch[0];
	wire [31:0] _r_T_5 = ~io_ea;
	wire _r_T_8 = io_bp_0_control_tmatch[0] & io_bp_0_address[0];
	wire _r_T_10 = (io_bp_0_control_tmatch[0] & io_bp_0_address[0]) & io_bp_0_address[1];
	wire _r_T_12 = ((io_bp_0_control_tmatch[0] & io_bp_0_address[0]) & io_bp_0_address[1]) & io_bp_0_address[2];
	wire [3:0] _r_T_13 = {_r_T_12, _r_T_10, _r_T_8, io_bp_0_control_tmatch[0]};
	wire [31:0] _GEN_11 = {28'd0, _r_T_13};
	wire [31:0] _r_T_14 = _r_T_5 | _GEN_11;
	wire [31:0] _r_T_15 = ~io_bp_0_address;
	wire [31:0] _r_T_24 = _r_T_15 | _GEN_11;
	wire _r_T_25 = _r_T_14 == _r_T_24;
	wire _r_T_26 = (io_bp_0_control_tmatch[1] ? _r_T_4 : _r_T_25);
	wire r = (en & io_bp_0_control_r) & _r_T_26;
	wire w = (en & io_bp_0_control_w) & _r_T_26;
	wire _x_T_4 = (io_pc >= io_bp_0_address) ^ io_bp_0_control_tmatch[0];
	wire [31:0] _x_T_5 = ~io_pc;
	wire [31:0] _x_T_14 = _x_T_5 | _GEN_11;
	wire _x_T_25 = _x_T_14 == _r_T_24;
	wire _x_T_26 = (io_bp_0_control_tmatch[1] ? _x_T_4 : _x_T_25);
	wire x = (en & io_bp_0_control_x) & _x_T_26;
	wire _io_xcpt_ld_T = ~io_bp_0_control_action;
	assign io_xcpt_if = x & _io_xcpt_ld_T;
	assign io_xcpt_ld = r & ~io_bp_0_control_action;
	assign io_xcpt_st = w & _io_xcpt_ld_T;
	assign io_debug_if = x & io_bp_0_control_action;
	assign io_debug_ld = r & io_bp_0_control_action;
	assign io_debug_st = w & io_bp_0_control_action;
endmodule
module ALU (
	io_fn,
	io_in2,
	io_in1,
	io_out,
	io_adder_out,
	io_cmp_out
);
	input [3:0] io_fn;
	input [31:0] io_in2;
	input [31:0] io_in1;
	output wire [31:0] io_out;
	output wire [31:0] io_adder_out;
	output wire io_cmp_out;
	wire [31:0] _in2_inv_T_1 = ~io_in2;
	wire [31:0] in2_inv = (io_fn[3] ? _in2_inv_T_1 : io_in2);
	wire [31:0] in1_xor_in2 = io_in1 ^ in2_inv;
	wire [31:0] _io_adder_out_T_1 = io_in1 + in2_inv;
	wire [31:0] _GEN_0 = {31'd0, io_fn[3]};
	wire _slt_T_7 = (io_fn[1] ? io_in2[31] : io_in1[31]);
	wire slt = (io_in1[31] == io_in2[31] ? io_adder_out[31] : _slt_T_7);
	wire _io_cmp_out_T_2 = ~io_fn[3];
	wire _io_cmp_out_T_4 = (_io_cmp_out_T_2 ? in1_xor_in2 == 32'h00000000 : slt);
	wire [4:0] shamt = io_in2[4:0];
	wire _shin_T_2 = (io_fn == 4'h5) | (io_fn == 4'hb);
	wire [31:0] _GEN_1 = {16'd0, io_in1[31:16]};
	wire [31:0] _shin_T_6 = _GEN_1 & 32'h0000ffff;
	wire [31:0] _shin_T_8 = {io_in1[15:0], 16'h0000};
	wire [31:0] _shin_T_10 = _shin_T_8 & 32'hffff0000;
	wire [31:0] _shin_T_11 = _shin_T_6 | _shin_T_10;
	wire [31:0] _GEN_2 = {8'd0, _shin_T_11[31:8]};
	wire [31:0] _shin_T_16 = _GEN_2 & 32'h00ff00ff;
	wire [31:0] _shin_T_18 = {_shin_T_11[23:0], 8'h00};
	wire [31:0] _shin_T_20 = _shin_T_18 & 32'hff00ff00;
	wire [31:0] _shin_T_21 = _shin_T_16 | _shin_T_20;
	wire [31:0] _GEN_3 = {4'd0, _shin_T_21[31:4]};
	wire [31:0] _shin_T_26 = _GEN_3 & 32'h0f0f0f0f;
	wire [31:0] _shin_T_28 = {_shin_T_21[27:0], 4'h0};
	wire [31:0] _shin_T_30 = _shin_T_28 & 32'hf0f0f0f0;
	wire [31:0] _shin_T_31 = _shin_T_26 | _shin_T_30;
	wire [31:0] _GEN_4 = {2'd0, _shin_T_31[31:2]};
	wire [31:0] _shin_T_36 = _GEN_4 & 32'h33333333;
	wire [31:0] _shin_T_38 = {_shin_T_31[29:0], 2'h0};
	wire [31:0] _shin_T_40 = _shin_T_38 & 32'hcccccccc;
	wire [31:0] _shin_T_41 = _shin_T_36 | _shin_T_40;
	wire [31:0] _GEN_5 = {1'd0, _shin_T_41[31:1]};
	wire [31:0] _shin_T_46 = _GEN_5 & 32'h55555555;
	wire [31:0] _shin_T_48 = {_shin_T_41[30:0], 1'h0};
	wire [31:0] _shin_T_50 = _shin_T_48 & 32'haaaaaaaa;
	wire [31:0] _shin_T_51 = _shin_T_46 | _shin_T_50;
	wire [31:0] shin = ((io_fn == 4'h5) | (io_fn == 4'hb) ? io_in1 : _shin_T_51);
	wire _shout_r_T_2 = io_fn[3] & shin[31];
	wire [32:0] _shout_r_T_4 = {_shout_r_T_2, shin};
	wire [32:0] _shout_r_T_5 = $signed(_shout_r_T_4) >>> shamt;
	wire [31:0] shout_r = _shout_r_T_5[31:0];
	wire [31:0] _GEN_6 = {16'd0, shout_r[31:16]};
	wire [31:0] _shout_l_T_3 = _GEN_6 & 32'h0000ffff;
	wire [31:0] _shout_l_T_5 = {shout_r[15:0], 16'h0000};
	wire [31:0] _shout_l_T_7 = _shout_l_T_5 & 32'hffff0000;
	wire [31:0] _shout_l_T_8 = _shout_l_T_3 | _shout_l_T_7;
	wire [31:0] _GEN_7 = {8'd0, _shout_l_T_8[31:8]};
	wire [31:0] _shout_l_T_13 = _GEN_7 & 32'h00ff00ff;
	wire [31:0] _shout_l_T_15 = {_shout_l_T_8[23:0], 8'h00};
	wire [31:0] _shout_l_T_17 = _shout_l_T_15 & 32'hff00ff00;
	wire [31:0] _shout_l_T_18 = _shout_l_T_13 | _shout_l_T_17;
	wire [31:0] _GEN_8 = {4'd0, _shout_l_T_18[31:4]};
	wire [31:0] _shout_l_T_23 = _GEN_8 & 32'h0f0f0f0f;
	wire [31:0] _shout_l_T_25 = {_shout_l_T_18[27:0], 4'h0};
	wire [31:0] _shout_l_T_27 = _shout_l_T_25 & 32'hf0f0f0f0;
	wire [31:0] _shout_l_T_28 = _shout_l_T_23 | _shout_l_T_27;
	wire [31:0] _GEN_9 = {2'd0, _shout_l_T_28[31:2]};
	wire [31:0] _shout_l_T_33 = _GEN_9 & 32'h33333333;
	wire [31:0] _shout_l_T_35 = {_shout_l_T_28[29:0], 2'h0};
	wire [31:0] _shout_l_T_37 = _shout_l_T_35 & 32'hcccccccc;
	wire [31:0] _shout_l_T_38 = _shout_l_T_33 | _shout_l_T_37;
	wire [31:0] _GEN_10 = {1'd0, _shout_l_T_38[31:1]};
	wire [31:0] _shout_l_T_43 = _GEN_10 & 32'h55555555;
	wire [31:0] _shout_l_T_45 = {_shout_l_T_38[30:0], 1'h0};
	wire [31:0] _shout_l_T_47 = _shout_l_T_45 & 32'haaaaaaaa;
	wire [31:0] shout_l = _shout_l_T_43 | _shout_l_T_47;
	wire [31:0] _shout_T_3 = (_shin_T_2 ? shout_r : 32'h00000000);
	wire [31:0] _shout_T_5 = (io_fn == 4'h1 ? shout_l : 32'h00000000);
	wire [31:0] shout = _shout_T_3 | _shout_T_5;
	wire _logic_T_1 = io_fn == 4'h6;
	wire [31:0] _logic_T_3 = ((io_fn == 4'h4) | (io_fn == 4'h6) ? in1_xor_in2 : 32'h00000000);
	wire [31:0] _logic_T_7 = io_in1 & io_in2;
	wire [31:0] _logic_T_8 = (_logic_T_1 | (io_fn == 4'h7) ? _logic_T_7 : 32'h00000000);
	wire [31:0] logic_ = _logic_T_3 | _logic_T_8;
	wire _shift_logic_T = io_fn >= 4'hc;
	wire _shift_logic_T_1 = _shift_logic_T & slt;
	wire [31:0] _GEN_11 = {31'd0, _shift_logic_T_1};
	wire [31:0] _shift_logic_T_2 = _GEN_11 | logic_;
	wire [31:0] shift_logic = _shift_logic_T_2 | shout;
	assign io_out = ((io_fn == 4'h0) | (io_fn == 4'ha) ? io_adder_out : shift_logic);
	assign io_adder_out = _io_adder_out_T_1 + _GEN_0;
	assign io_cmp_out = io_fn[0] ^ _io_cmp_out_T_4;
endmodule
module MulDiv (
	clock,
	reset,
	io_req_ready,
	io_req_valid,
	io_req_bits_fn,
	io_req_bits_in1,
	io_req_bits_in2,
	io_req_bits_tag,
	io_kill,
	io_resp_ready,
	io_resp_valid,
	io_resp_bits_data,
	io_resp_bits_tag
);
	input clock;
	input reset;
	output wire io_req_ready;
	input io_req_valid;
	input [3:0] io_req_bits_fn;
	input [31:0] io_req_bits_in1;
	input [31:0] io_req_bits_in2;
	input [4:0] io_req_bits_tag;
	input io_kill;
	input io_resp_ready;
	output wire io_resp_valid;
	output wire [31:0] io_resp_bits_data;
	output wire [4:0] io_resp_bits_tag;
	reg [2:0] state;
	reg [4:0] req_tag;
	reg [5:0] count;
	reg neg_out;
	reg isHi;
	reg resHi;
	reg [32:0] divisor;
	reg [65:0] remainder;
	wire [3:0] _T = io_req_bits_fn & 4'h4;
	wire cmdMul = _T == 4'h0;
	wire [3:0] _T_3 = io_req_bits_fn & 4'h5;
	wire _T_4 = _T_3 == 4'h1;
	wire [3:0] _T_5 = io_req_bits_fn & 4'h2;
	wire _T_6 = _T_5 == 4'h2;
	wire cmdHi = _T_4 | _T_6;
	wire [3:0] _T_9 = io_req_bits_fn & 4'h6;
	wire _T_10 = _T_9 == 4'h0;
	wire [3:0] _T_11 = io_req_bits_fn & 4'h1;
	wire _T_12 = _T_11 == 4'h0;
	wire lhsSigned = _T_10 | _T_12;
	wire _T_16 = _T_3 == 4'h4;
	wire rhsSigned = _T_10 | _T_16;
	wire lhs_sign = lhsSigned & io_req_bits_in1[31];
	wire [15:0] hi = io_req_bits_in1[31:16];
	wire [31:0] lhs_in = {hi, io_req_bits_in1[15:0]};
	wire rhs_sign = rhsSigned & io_req_bits_in2[31];
	wire [15:0] hi_1 = io_req_bits_in2[31:16];
	wire [32:0] subtractor = remainder[64:32] - divisor;
	wire [31:0] result = (resHi ? remainder[64:33] : remainder[31:0]);
	wire [31:0] negated_remainder = 32'h00000000 - result;
	wire [65:0] _GEN_0 = (remainder[31] ? {34'd0, negated_remainder} : remainder);
	wire [65:0] _GEN_2 = (state == 3'h1 ? _GEN_0 : remainder);
	wire [2:0] _GEN_4 = (state == 3'h1 ? 3'h3 : state);
	wire [2:0] _GEN_6 = (state == 3'h5 ? 3'h7 : _GEN_4);
	wire _GEN_7 = (state == 3'h5 ? 1'h0 : resHi);
	wire [64:0] mulReg = {remainder[65:33], remainder[31:0]};
	wire mplierSign = remainder[32];
	wire [31:0] mplier = mulReg[31:0];
	wire [32:0] accum = mulReg[64:32];
	wire [8:0] _prod_T_2 = {mplierSign, mplier[7:0]};
	wire [41:0] _prod_T_3 = $signed(_prod_T_2) * $signed(divisor);
	wire [41:0] _GEN_35 = {{9 {accum[32]}}, accum};
	wire [41:0] nextMulReg_hi = $signed(_prod_T_3) + $signed(_GEN_35);
	wire [65:0] nextMulReg = {nextMulReg_hi, mplier[31:8]};
	wire nextMplierSign = (count == 6'h02) & neg_out;
	wire _eOut_T_4 = ~isHi;
	wire [64:0] nextMulReg1 = {nextMulReg[64:32], nextMulReg[31:0]};
	wire [65:0] _remainder_T_2 = {nextMulReg1[64:32], nextMplierSign, nextMulReg1[31:0]};
	wire [5:0] _count_T_1 = count + 6'h01;
	wire [2:0] _GEN_8 = (count == 6'h03 ? 3'h6 : _GEN_6);
	wire _GEN_9 = (count == 6'h03 ? isHi : _GEN_7);
	wire [2:0] _GEN_12 = (state == 3'h2 ? _GEN_8 : _GEN_6);
	wire _GEN_13 = (state == 3'h2 ? _GEN_9 : _GEN_7);
	wire unrolls_less = subtractor[32];
	wire [31:0] _unrolls_T_2 = (unrolls_less ? remainder[63:32] : subtractor[31:0]);
	wire _unrolls_T_4 = ~unrolls_less;
	wire [64:0] unrolls_0 = {_unrolls_T_2, remainder[31:0], _unrolls_T_4};
	wire [2:0] _state_T = (neg_out ? 3'h5 : 3'h7);
	wire [2:0] _GEN_14 = (count == 6'h20 ? _state_T : _GEN_12);
	wire divby0 = (count == 6'h00) & _unrolls_T_4;
	wire _T_36 = io_resp_ready & io_resp_valid;
	wire _T_38 = io_req_ready & io_req_valid;
	wire [32:0] _divisor_T = {rhs_sign, hi_1, io_req_bits_in2[15:0]};
	wire [15:0] loOut = result[15:0];
	assign io_req_ready = state == 3'h0;
	assign io_resp_valid = (state == 3'h6) | (state == 3'h7);
	assign io_resp_bits_data = {result[31:16], loOut};
	assign io_resp_bits_tag = req_tag;
	always @(posedge clock) begin
		if (reset)
			state <= 3'h0;
		else if (_T_38) begin
			if (cmdMul)
				state <= 3'h2;
			else if (lhs_sign | rhs_sign)
				state <= 3'h1;
			else
				state <= 3'h3;
		end
		else if (_T_36 | io_kill)
			state <= 3'h0;
		else if (state == 3'h3)
			state <= _GEN_14;
		else
			state <= _GEN_12;
		if (_T_38)
			req_tag <= io_req_bits_tag;
		if (_T_38)
			count <= 6'h00;
		else if (state == 3'h3)
			count <= _count_T_1;
		else if (state == 3'h2)
			count <= _count_T_1;
		if (_T_38) begin
			if (cmdHi)
				neg_out <= lhs_sign;
			else
				neg_out <= lhs_sign != rhs_sign;
		end
		else if (state == 3'h3)
			if (divby0 & _eOut_T_4)
				neg_out <= 1'h0;
		if (_T_38)
			isHi <= cmdHi;
		if (_T_38)
			resHi <= 1'h0;
		else if (state == 3'h3) begin
			if (count == 6'h20)
				resHi <= isHi;
			else
				resHi <= _GEN_13;
		end
		else
			resHi <= _GEN_13;
		if (_T_38)
			divisor <= _divisor_T;
		else if (state == 3'h1)
			if (divisor[31])
				divisor <= subtractor;
		if (_T_38)
			remainder <= {34'd0, lhs_in};
		else if (state == 3'h3)
			remainder <= {1'd0, unrolls_0};
		else if (state == 3'h2)
			remainder <= _remainder_T_2;
		else if (state == 3'h5)
			remainder <= {34'd0, negated_remainder};
		else
			remainder <= _GEN_2;
	end
endmodule
module PlusArgTimeout (
	clock,
	reset,
	io_count
);
	input clock;
	input reset;
	input [31:0] io_count;
	wire [31:0] plusarg_reader_out;
	wire _T = plusarg_reader_out > 32'h00000000;
	plusarg_reader #(
		.FORMAT("max_core_cycles=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	always @(posedge clock)
		;
endmodule
module Rocket (
	clock,
	reset,
	io_hartid,
	io_interrupts_debug,
	io_interrupts_mtip,
	io_interrupts_msip,
	io_interrupts_meip,
	io_imem_might_request,
	io_imem_req_valid,
	io_imem_req_bits_pc,
	io_imem_req_bits_speculative,
	io_imem_resp_ready,
	io_imem_resp_valid,
	io_imem_resp_bits_pc,
	io_imem_resp_bits_data,
	io_imem_resp_bits_xcpt_ae_inst,
	io_imem_resp_bits_replay,
	io_imem_btb_update_valid,
	io_imem_bht_update_valid,
	io_imem_flush_icache,
	io_dmem_req_ready,
	io_dmem_req_valid,
	io_dmem_req_bits_addr,
	io_dmem_req_bits_tag,
	io_dmem_req_bits_cmd,
	io_dmem_req_bits_size,
	io_dmem_req_bits_signed,
	io_dmem_req_bits_dv,
	io_dmem_s1_kill,
	io_dmem_s1_data_data,
	io_dmem_s2_nack,
	io_dmem_resp_valid,
	io_dmem_resp_bits_tag,
	io_dmem_resp_bits_data,
	io_dmem_resp_bits_replay,
	io_dmem_resp_bits_has_data,
	io_dmem_resp_bits_data_word_bypass,
	io_dmem_replay_next,
	io_dmem_s2_xcpt_ma_ld,
	io_dmem_s2_xcpt_ma_st,
	io_dmem_s2_xcpt_pf_ld,
	io_dmem_s2_xcpt_pf_st,
	io_dmem_s2_xcpt_ae_ld,
	io_dmem_s2_xcpt_ae_st,
	io_dmem_ordered,
	io_dmem_perf_grant,
	io_ptw_status_debug,
	io_ptw_pmp_0_cfg_l,
	io_ptw_pmp_0_cfg_a,
	io_ptw_pmp_0_cfg_x,
	io_ptw_pmp_0_cfg_w,
	io_ptw_pmp_0_cfg_r,
	io_ptw_pmp_0_addr,
	io_ptw_pmp_0_mask,
	io_ptw_pmp_1_cfg_l,
	io_ptw_pmp_1_cfg_a,
	io_ptw_pmp_1_cfg_x,
	io_ptw_pmp_1_cfg_w,
	io_ptw_pmp_1_cfg_r,
	io_ptw_pmp_1_addr,
	io_ptw_pmp_1_mask,
	io_ptw_pmp_2_cfg_l,
	io_ptw_pmp_2_cfg_a,
	io_ptw_pmp_2_cfg_x,
	io_ptw_pmp_2_cfg_w,
	io_ptw_pmp_2_cfg_r,
	io_ptw_pmp_2_addr,
	io_ptw_pmp_2_mask,
	io_ptw_pmp_3_cfg_l,
	io_ptw_pmp_3_cfg_a,
	io_ptw_pmp_3_cfg_x,
	io_ptw_pmp_3_cfg_w,
	io_ptw_pmp_3_cfg_r,
	io_ptw_pmp_3_addr,
	io_ptw_pmp_3_mask,
	io_ptw_pmp_4_cfg_l,
	io_ptw_pmp_4_cfg_a,
	io_ptw_pmp_4_cfg_x,
	io_ptw_pmp_4_cfg_w,
	io_ptw_pmp_4_cfg_r,
	io_ptw_pmp_4_addr,
	io_ptw_pmp_4_mask,
	io_ptw_pmp_5_cfg_l,
	io_ptw_pmp_5_cfg_a,
	io_ptw_pmp_5_cfg_x,
	io_ptw_pmp_5_cfg_w,
	io_ptw_pmp_5_cfg_r,
	io_ptw_pmp_5_addr,
	io_ptw_pmp_5_mask,
	io_ptw_pmp_6_cfg_l,
	io_ptw_pmp_6_cfg_a,
	io_ptw_pmp_6_cfg_x,
	io_ptw_pmp_6_cfg_w,
	io_ptw_pmp_6_cfg_r,
	io_ptw_pmp_6_addr,
	io_ptw_pmp_6_mask,
	io_ptw_pmp_7_cfg_l,
	io_ptw_pmp_7_cfg_a,
	io_ptw_pmp_7_cfg_x,
	io_ptw_pmp_7_cfg_w,
	io_ptw_pmp_7_cfg_r,
	io_ptw_pmp_7_addr,
	io_ptw_pmp_7_mask,
	io_ptw_customCSRs_csrs_0_value,
	io_wfi
);
	input clock;
	input reset;
	input io_hartid;
	input io_interrupts_debug;
	input io_interrupts_mtip;
	input io_interrupts_msip;
	input io_interrupts_meip;
	output wire io_imem_might_request;
	output wire io_imem_req_valid;
	output wire [31:0] io_imem_req_bits_pc;
	output wire io_imem_req_bits_speculative;
	output wire io_imem_resp_ready;
	input io_imem_resp_valid;
	input [31:0] io_imem_resp_bits_pc;
	input [31:0] io_imem_resp_bits_data;
	input io_imem_resp_bits_xcpt_ae_inst;
	input io_imem_resp_bits_replay;
	output wire io_imem_btb_update_valid;
	output wire io_imem_bht_update_valid;
	output wire io_imem_flush_icache;
	input io_dmem_req_ready;
	output wire io_dmem_req_valid;
	output wire [31:0] io_dmem_req_bits_addr;
	output wire [6:0] io_dmem_req_bits_tag;
	output wire [4:0] io_dmem_req_bits_cmd;
	output wire [1:0] io_dmem_req_bits_size;
	output wire io_dmem_req_bits_signed;
	output wire io_dmem_req_bits_dv;
	output wire io_dmem_s1_kill;
	output wire [31:0] io_dmem_s1_data_data;
	input io_dmem_s2_nack;
	input io_dmem_resp_valid;
	input [6:0] io_dmem_resp_bits_tag;
	input [31:0] io_dmem_resp_bits_data;
	input io_dmem_resp_bits_replay;
	input io_dmem_resp_bits_has_data;
	input [31:0] io_dmem_resp_bits_data_word_bypass;
	input io_dmem_replay_next;
	input io_dmem_s2_xcpt_ma_ld;
	input io_dmem_s2_xcpt_ma_st;
	input io_dmem_s2_xcpt_pf_ld;
	input io_dmem_s2_xcpt_pf_st;
	input io_dmem_s2_xcpt_ae_ld;
	input io_dmem_s2_xcpt_ae_st;
	input io_dmem_ordered;
	input io_dmem_perf_grant;
	output wire io_ptw_status_debug;
	output wire io_ptw_pmp_0_cfg_l;
	output wire [1:0] io_ptw_pmp_0_cfg_a;
	output wire io_ptw_pmp_0_cfg_x;
	output wire io_ptw_pmp_0_cfg_w;
	output wire io_ptw_pmp_0_cfg_r;
	output wire [29:0] io_ptw_pmp_0_addr;
	output wire [31:0] io_ptw_pmp_0_mask;
	output wire io_ptw_pmp_1_cfg_l;
	output wire [1:0] io_ptw_pmp_1_cfg_a;
	output wire io_ptw_pmp_1_cfg_x;
	output wire io_ptw_pmp_1_cfg_w;
	output wire io_ptw_pmp_1_cfg_r;
	output wire [29:0] io_ptw_pmp_1_addr;
	output wire [31:0] io_ptw_pmp_1_mask;
	output wire io_ptw_pmp_2_cfg_l;
	output wire [1:0] io_ptw_pmp_2_cfg_a;
	output wire io_ptw_pmp_2_cfg_x;
	output wire io_ptw_pmp_2_cfg_w;
	output wire io_ptw_pmp_2_cfg_r;
	output wire [29:0] io_ptw_pmp_2_addr;
	output wire [31:0] io_ptw_pmp_2_mask;
	output wire io_ptw_pmp_3_cfg_l;
	output wire [1:0] io_ptw_pmp_3_cfg_a;
	output wire io_ptw_pmp_3_cfg_x;
	output wire io_ptw_pmp_3_cfg_w;
	output wire io_ptw_pmp_3_cfg_r;
	output wire [29:0] io_ptw_pmp_3_addr;
	output wire [31:0] io_ptw_pmp_3_mask;
	output wire io_ptw_pmp_4_cfg_l;
	output wire [1:0] io_ptw_pmp_4_cfg_a;
	output wire io_ptw_pmp_4_cfg_x;
	output wire io_ptw_pmp_4_cfg_w;
	output wire io_ptw_pmp_4_cfg_r;
	output wire [29:0] io_ptw_pmp_4_addr;
	output wire [31:0] io_ptw_pmp_4_mask;
	output wire io_ptw_pmp_5_cfg_l;
	output wire [1:0] io_ptw_pmp_5_cfg_a;
	output wire io_ptw_pmp_5_cfg_x;
	output wire io_ptw_pmp_5_cfg_w;
	output wire io_ptw_pmp_5_cfg_r;
	output wire [29:0] io_ptw_pmp_5_addr;
	output wire [31:0] io_ptw_pmp_5_mask;
	output wire io_ptw_pmp_6_cfg_l;
	output wire [1:0] io_ptw_pmp_6_cfg_a;
	output wire io_ptw_pmp_6_cfg_x;
	output wire io_ptw_pmp_6_cfg_w;
	output wire io_ptw_pmp_6_cfg_r;
	output wire [29:0] io_ptw_pmp_6_addr;
	output wire [31:0] io_ptw_pmp_6_mask;
	output wire io_ptw_pmp_7_cfg_l;
	output wire [1:0] io_ptw_pmp_7_cfg_a;
	output wire io_ptw_pmp_7_cfg_x;
	output wire io_ptw_pmp_7_cfg_w;
	output wire io_ptw_pmp_7_cfg_r;
	output wire [29:0] io_ptw_pmp_7_addr;
	output wire [31:0] io_ptw_pmp_7_mask;
	output wire [31:0] io_ptw_customCSRs_csrs_0_value;
	output wire io_wfi;
	wire ibuf_clock;
	wire ibuf_reset;
	wire ibuf_io_imem_ready;
	wire ibuf_io_imem_valid;
	wire [31:0] ibuf_io_imem_bits_pc;
	wire [31:0] ibuf_io_imem_bits_data;
	wire ibuf_io_imem_bits_xcpt_ae_inst;
	wire ibuf_io_imem_bits_replay;
	wire ibuf_io_kill;
	wire [31:0] ibuf_io_pc;
	wire ibuf_io_inst_0_ready;
	wire ibuf_io_inst_0_valid;
	wire ibuf_io_inst_0_bits_xcpt0_ae_inst;
	wire ibuf_io_inst_0_bits_xcpt1_pf_inst;
	wire ibuf_io_inst_0_bits_xcpt1_gf_inst;
	wire ibuf_io_inst_0_bits_xcpt1_ae_inst;
	wire ibuf_io_inst_0_bits_replay;
	wire ibuf_io_inst_0_bits_rvc;
	wire [31:0] ibuf_io_inst_0_bits_inst_bits;
	wire [4:0] ibuf_io_inst_0_bits_inst_rd;
	wire [4:0] ibuf_io_inst_0_bits_inst_rs1;
	wire [4:0] ibuf_io_inst_0_bits_inst_rs2;
	wire [31:0] ibuf_io_inst_0_bits_raw;
	reg [31:0] rf [0:30];
	wire rf_id_rs_MPORT_en;
	wire [4:0] rf_id_rs_MPORT_addr;
	wire [31:0] rf_id_rs_MPORT_data;
	wire rf_id_rs_MPORT_1_en;
	wire [4:0] rf_id_rs_MPORT_1_addr;
	wire [31:0] rf_id_rs_MPORT_1_data;
	wire [31:0] rf_MPORT_data;
	wire [4:0] rf_MPORT_addr;
	wire rf_MPORT_mask;
	wire rf_MPORT_en;
	wire csr_clock;
	wire csr_reset;
	wire csr_io_ungated_clock;
	wire csr_io_interrupts_debug;
	wire csr_io_interrupts_mtip;
	wire csr_io_interrupts_msip;
	wire csr_io_interrupts_meip;
	wire csr_io_hartid;
	wire [11:0] csr_io_rw_addr;
	wire [2:0] csr_io_rw_cmd;
	wire [31:0] csr_io_rw_rdata;
	wire [31:0] csr_io_rw_wdata;
	wire [31:0] csr_io_decode_0_inst;
	wire csr_io_decode_0_fp_illegal;
	wire csr_io_decode_0_fp_csr;
	wire csr_io_decode_0_read_illegal;
	wire csr_io_decode_0_write_illegal;
	wire csr_io_decode_0_write_flush;
	wire csr_io_decode_0_system_illegal;
	wire csr_io_csr_stall;
	wire csr_io_eret;
	wire csr_io_singleStep;
	wire csr_io_status_debug;
	wire csr_io_status_cease;
	wire csr_io_status_wfi;
	wire [31:0] csr_io_status_isa;
	wire [1:0] csr_io_status_dprv;
	wire csr_io_status_dv;
	wire [1:0] csr_io_status_prv;
	wire csr_io_status_v;
	wire csr_io_status_sd;
	wire [22:0] csr_io_status_zero2;
	wire csr_io_status_mpv;
	wire csr_io_status_gva;
	wire csr_io_status_mbe;
	wire csr_io_status_sbe;
	wire [1:0] csr_io_status_sxl;
	wire [1:0] csr_io_status_uxl;
	wire csr_io_status_sd_rv32;
	wire [7:0] csr_io_status_zero1;
	wire csr_io_status_tsr;
	wire csr_io_status_tw;
	wire csr_io_status_tvm;
	wire csr_io_status_mxr;
	wire csr_io_status_sum;
	wire csr_io_status_mprv;
	wire [1:0] csr_io_status_xs;
	wire [1:0] csr_io_status_fs;
	wire [1:0] csr_io_status_mpp;
	wire [1:0] csr_io_status_vs;
	wire csr_io_status_spp;
	wire csr_io_status_mpie;
	wire csr_io_status_ube;
	wire csr_io_status_spie;
	wire csr_io_status_upie;
	wire csr_io_status_mie;
	wire csr_io_status_hie;
	wire csr_io_status_sie;
	wire csr_io_status_uie;
	wire [31:0] csr_io_evec;
	wire csr_io_exception;
	wire csr_io_retire;
	wire [31:0] csr_io_cause;
	wire [31:0] csr_io_pc;
	wire [31:0] csr_io_tval;
	wire csr_io_gva;
	wire [31:0] csr_io_time;
	wire csr_io_interrupt;
	wire [31:0] csr_io_interrupt_cause;
	wire csr_io_bp_0_control_action;
	wire [1:0] csr_io_bp_0_control_tmatch;
	wire csr_io_bp_0_control_x;
	wire csr_io_bp_0_control_w;
	wire csr_io_bp_0_control_r;
	wire [31:0] csr_io_bp_0_address;
	wire csr_io_pmp_0_cfg_l;
	wire [1:0] csr_io_pmp_0_cfg_a;
	wire csr_io_pmp_0_cfg_x;
	wire csr_io_pmp_0_cfg_w;
	wire csr_io_pmp_0_cfg_r;
	wire [29:0] csr_io_pmp_0_addr;
	wire [31:0] csr_io_pmp_0_mask;
	wire csr_io_pmp_1_cfg_l;
	wire [1:0] csr_io_pmp_1_cfg_a;
	wire csr_io_pmp_1_cfg_x;
	wire csr_io_pmp_1_cfg_w;
	wire csr_io_pmp_1_cfg_r;
	wire [29:0] csr_io_pmp_1_addr;
	wire [31:0] csr_io_pmp_1_mask;
	wire csr_io_pmp_2_cfg_l;
	wire [1:0] csr_io_pmp_2_cfg_a;
	wire csr_io_pmp_2_cfg_x;
	wire csr_io_pmp_2_cfg_w;
	wire csr_io_pmp_2_cfg_r;
	wire [29:0] csr_io_pmp_2_addr;
	wire [31:0] csr_io_pmp_2_mask;
	wire csr_io_pmp_3_cfg_l;
	wire [1:0] csr_io_pmp_3_cfg_a;
	wire csr_io_pmp_3_cfg_x;
	wire csr_io_pmp_3_cfg_w;
	wire csr_io_pmp_3_cfg_r;
	wire [29:0] csr_io_pmp_3_addr;
	wire [31:0] csr_io_pmp_3_mask;
	wire csr_io_pmp_4_cfg_l;
	wire [1:0] csr_io_pmp_4_cfg_a;
	wire csr_io_pmp_4_cfg_x;
	wire csr_io_pmp_4_cfg_w;
	wire csr_io_pmp_4_cfg_r;
	wire [29:0] csr_io_pmp_4_addr;
	wire [31:0] csr_io_pmp_4_mask;
	wire csr_io_pmp_5_cfg_l;
	wire [1:0] csr_io_pmp_5_cfg_a;
	wire csr_io_pmp_5_cfg_x;
	wire csr_io_pmp_5_cfg_w;
	wire csr_io_pmp_5_cfg_r;
	wire [29:0] csr_io_pmp_5_addr;
	wire [31:0] csr_io_pmp_5_mask;
	wire csr_io_pmp_6_cfg_l;
	wire [1:0] csr_io_pmp_6_cfg_a;
	wire csr_io_pmp_6_cfg_x;
	wire csr_io_pmp_6_cfg_w;
	wire csr_io_pmp_6_cfg_r;
	wire [29:0] csr_io_pmp_6_addr;
	wire [31:0] csr_io_pmp_6_mask;
	wire csr_io_pmp_7_cfg_l;
	wire [1:0] csr_io_pmp_7_cfg_a;
	wire csr_io_pmp_7_cfg_x;
	wire csr_io_pmp_7_cfg_w;
	wire csr_io_pmp_7_cfg_r;
	wire [29:0] csr_io_pmp_7_addr;
	wire [31:0] csr_io_pmp_7_mask;
	wire csr_io_inhibit_cycle;
	wire [31:0] csr_io_inst_0;
	wire csr_io_trace_0_valid;
	wire [31:0] csr_io_trace_0_iaddr;
	wire [31:0] csr_io_trace_0_insn;
	wire csr_io_trace_0_exception;
	wire [31:0] csr_io_customCSRs_0_value;
	wire bpu_io_status_debug;
	wire bpu_io_bp_0_control_action;
	wire [1:0] bpu_io_bp_0_control_tmatch;
	wire bpu_io_bp_0_control_x;
	wire bpu_io_bp_0_control_w;
	wire bpu_io_bp_0_control_r;
	wire [31:0] bpu_io_bp_0_address;
	wire [31:0] bpu_io_pc;
	wire [31:0] bpu_io_ea;
	wire bpu_io_xcpt_if;
	wire bpu_io_xcpt_ld;
	wire bpu_io_xcpt_st;
	wire bpu_io_debug_if;
	wire bpu_io_debug_ld;
	wire bpu_io_debug_st;
	wire [3:0] alu_io_fn;
	wire [31:0] alu_io_in2;
	wire [31:0] alu_io_in1;
	wire [31:0] alu_io_out;
	wire [31:0] alu_io_adder_out;
	wire alu_io_cmp_out;
	wire div_clock;
	wire div_reset;
	wire div_io_req_ready;
	wire div_io_req_valid;
	wire [3:0] div_io_req_bits_fn;
	wire [31:0] div_io_req_bits_in1;
	wire [31:0] div_io_req_bits_in2;
	wire [4:0] div_io_req_bits_tag;
	wire div_io_kill;
	wire div_io_resp_ready;
	wire div_io_resp_valid;
	wire [31:0] div_io_resp_bits_data;
	wire [4:0] div_io_resp_bits_tag;
	wire PlusArgTimeout_clock;
	wire PlusArgTimeout_reset;
	wire [31:0] PlusArgTimeout_io_count;
	reg id_reg_pause;
	reg imem_might_request_reg;
	reg ex_ctrl_branch;
	reg ex_ctrl_jal;
	reg ex_ctrl_jalr;
	reg ex_ctrl_rxs2;
	reg ex_ctrl_rxs1;
	reg [1:0] ex_ctrl_sel_alu2;
	reg [1:0] ex_ctrl_sel_alu1;
	reg [2:0] ex_ctrl_sel_imm;
	reg [3:0] ex_ctrl_alu_fn;
	reg ex_ctrl_mem;
	reg [4:0] ex_ctrl_mem_cmd;
	reg ex_ctrl_div;
	reg ex_ctrl_wxd;
	reg [2:0] ex_ctrl_csr;
	reg ex_ctrl_fence_i;
	reg mem_ctrl_branch;
	reg mem_ctrl_jal;
	reg mem_ctrl_jalr;
	reg mem_ctrl_rxs2;
	reg mem_ctrl_rxs1;
	reg mem_ctrl_mem;
	reg mem_ctrl_div;
	reg mem_ctrl_wxd;
	reg [2:0] mem_ctrl_csr;
	reg mem_ctrl_fence_i;
	reg wb_ctrl_rxs2;
	reg wb_ctrl_rxs1;
	reg wb_ctrl_mem;
	reg wb_ctrl_div;
	reg wb_ctrl_wxd;
	reg [2:0] wb_ctrl_csr;
	reg wb_ctrl_fence_i;
	reg ex_reg_xcpt_interrupt;
	reg ex_reg_valid;
	reg ex_reg_rvc;
	reg ex_reg_xcpt;
	reg ex_reg_flush_pipe;
	reg ex_reg_load_use;
	reg [31:0] ex_reg_cause;
	reg ex_reg_replay;
	reg [31:0] ex_reg_pc;
	reg [1:0] ex_reg_mem_size;
	reg [31:0] ex_reg_inst;
	reg [31:0] ex_reg_raw_inst;
	reg mem_reg_xcpt_interrupt;
	reg mem_reg_valid;
	reg mem_reg_rvc;
	reg mem_reg_xcpt;
	reg mem_reg_replay;
	reg mem_reg_flush_pipe;
	reg [31:0] mem_reg_cause;
	reg mem_reg_slow_bypass;
	reg mem_reg_load;
	reg mem_reg_store;
	reg [31:0] mem_reg_pc;
	reg [31:0] mem_reg_inst;
	reg mem_reg_hls_or_dv;
	reg [31:0] mem_reg_raw_inst;
	reg [31:0] mem_reg_wdata;
	reg [31:0] mem_reg_rs2;
	reg mem_br_taken;
	reg wb_reg_valid;
	reg wb_reg_xcpt;
	reg wb_reg_replay;
	reg wb_reg_flush_pipe;
	reg [31:0] wb_reg_cause;
	reg [31:0] wb_reg_pc;
	reg wb_reg_hls_or_dv;
	reg [31:0] wb_reg_inst;
	reg [31:0] wb_reg_raw_inst;
	reg [31:0] wb_reg_wdata;
	wire replay_wb_common = io_dmem_s2_nack | wb_reg_replay;
	wire _T_90 = wb_reg_valid & wb_ctrl_mem;
	wire _T_91 = (wb_reg_valid & wb_ctrl_mem) & io_dmem_s2_xcpt_pf_st;
	wire _T_93 = _T_90 & io_dmem_s2_xcpt_pf_ld;
	wire _T_99 = _T_90 & io_dmem_s2_xcpt_ae_st;
	wire _T_101 = _T_90 & io_dmem_s2_xcpt_ae_ld;
	wire _T_103 = _T_90 & io_dmem_s2_xcpt_ma_st;
	wire _T_105 = _T_90 & io_dmem_s2_xcpt_ma_ld;
	wire wb_xcpt = (((((wb_reg_xcpt | _T_91) | _T_93) | _T_99) | _T_101) | _T_103) | _T_105;
	wire take_pc_wb = ((replay_wb_common | wb_xcpt) | csr_io_eret) | wb_reg_flush_pipe;
	wire _take_pc_mem_T = ~mem_reg_xcpt;
	wire _mem_cfi_taken_T = mem_ctrl_branch & mem_br_taken;
	wire mem_cfi_taken = ((mem_ctrl_branch & mem_br_taken) | mem_ctrl_jalr) | mem_ctrl_jal;
	wire take_pc_mem = (mem_reg_valid & ~mem_reg_xcpt) & mem_cfi_taken;
	wire take_pc_mem_wb = take_pc_wb | take_pc_mem;
	wire [31:0] _id_ctrl_decoder_bit_T = ibuf_io_inst_0_bits_inst_bits & 32'hfe00707f;
	wire _id_ctrl_decoder_bit_T_1 = _id_ctrl_decoder_bit_T == 32'h02000033;
	wire _id_ctrl_decoder_bit_T_3 = _id_ctrl_decoder_bit_T == 32'h02001033;
	wire _id_ctrl_decoder_bit_T_5 = _id_ctrl_decoder_bit_T == 32'h02003033;
	wire _id_ctrl_decoder_bit_T_7 = _id_ctrl_decoder_bit_T == 32'h02002033;
	wire _id_ctrl_decoder_bit_T_9 = _id_ctrl_decoder_bit_T == 32'h02004033;
	wire _id_ctrl_decoder_bit_T_11 = _id_ctrl_decoder_bit_T == 32'h02005033;
	wire _id_ctrl_decoder_bit_T_13 = _id_ctrl_decoder_bit_T == 32'h02006033;
	wire _id_ctrl_decoder_bit_T_15 = _id_ctrl_decoder_bit_T == 32'h02007033;
	wire [31:0] _id_ctrl_decoder_bit_T_16 = ibuf_io_inst_0_bits_inst_bits & 32'hf800707f;
	wire _id_ctrl_decoder_bit_T_17 = _id_ctrl_decoder_bit_T_16 == 32'h0000202f;
	wire _id_ctrl_decoder_bit_T_19 = _id_ctrl_decoder_bit_T_16 == 32'h2000202f;
	wire _id_ctrl_decoder_bit_T_21 = _id_ctrl_decoder_bit_T_16 == 32'h0800202f;
	wire _id_ctrl_decoder_bit_T_23 = _id_ctrl_decoder_bit_T_16 == 32'h6000202f;
	wire _id_ctrl_decoder_bit_T_25 = _id_ctrl_decoder_bit_T_16 == 32'h4000202f;
	wire _id_ctrl_decoder_bit_T_27 = _id_ctrl_decoder_bit_T_16 == 32'h8000202f;
	wire _id_ctrl_decoder_bit_T_29 = _id_ctrl_decoder_bit_T_16 == 32'hc000202f;
	wire _id_ctrl_decoder_bit_T_31 = _id_ctrl_decoder_bit_T_16 == 32'ha000202f;
	wire _id_ctrl_decoder_bit_T_33 = _id_ctrl_decoder_bit_T_16 == 32'he000202f;
	wire [31:0] _id_ctrl_decoder_bit_T_34 = ibuf_io_inst_0_bits_inst_bits & 32'hf9f0707f;
	wire _id_ctrl_decoder_bit_T_35 = _id_ctrl_decoder_bit_T_34 == 32'h1000202f;
	wire _id_ctrl_decoder_bit_T_37 = _id_ctrl_decoder_bit_T_16 == 32'h1800202f;
	wire _id_ctrl_decoder_bit_T_39 = _id_ctrl_decoder_bit_T == 32'h00001013;
	wire _id_ctrl_decoder_bit_T_41 = _id_ctrl_decoder_bit_T == 32'h00005013;
	wire _id_ctrl_decoder_bit_T_43 = _id_ctrl_decoder_bit_T == 32'h40005013;
	wire _id_ctrl_decoder_bit_T_44 = ibuf_io_inst_0_bits_inst_bits == 32'h7b200073;
	wire [31:0] _id_ctrl_decoder_bit_T_45 = ibuf_io_inst_0_bits_inst_bits & 32'h0000707f;
	wire _id_ctrl_decoder_bit_T_46 = _id_ctrl_decoder_bit_T_45 == 32'h0000100f;
	wire _id_ctrl_decoder_bit_T_48 = _id_ctrl_decoder_bit_T_45 == 32'h00001063;
	wire _id_ctrl_decoder_bit_T_50 = _id_ctrl_decoder_bit_T_45 == 32'h00000063;
	wire _id_ctrl_decoder_bit_T_52 = _id_ctrl_decoder_bit_T_45 == 32'h00004063;
	wire _id_ctrl_decoder_bit_T_54 = _id_ctrl_decoder_bit_T_45 == 32'h00006063;
	wire _id_ctrl_decoder_bit_T_56 = _id_ctrl_decoder_bit_T_45 == 32'h00005063;
	wire _id_ctrl_decoder_bit_T_58 = _id_ctrl_decoder_bit_T_45 == 32'h00007063;
	wire [31:0] _id_ctrl_decoder_bit_T_59 = ibuf_io_inst_0_bits_inst_bits & 32'h0000007f;
	wire _id_ctrl_decoder_bit_T_60 = _id_ctrl_decoder_bit_T_59 == 32'h0000006f;
	wire _id_ctrl_decoder_bit_T_62 = _id_ctrl_decoder_bit_T_45 == 32'h00000067;
	wire _id_ctrl_decoder_bit_T_64 = _id_ctrl_decoder_bit_T_59 == 32'h00000017;
	wire _id_ctrl_decoder_bit_T_66 = _id_ctrl_decoder_bit_T_45 == 32'h00000003;
	wire _id_ctrl_decoder_bit_T_68 = _id_ctrl_decoder_bit_T_45 == 32'h00001003;
	wire _id_ctrl_decoder_bit_T_70 = _id_ctrl_decoder_bit_T_45 == 32'h00002003;
	wire _id_ctrl_decoder_bit_T_72 = _id_ctrl_decoder_bit_T_45 == 32'h00004003;
	wire _id_ctrl_decoder_bit_T_74 = _id_ctrl_decoder_bit_T_45 == 32'h00005003;
	wire _id_ctrl_decoder_bit_T_76 = _id_ctrl_decoder_bit_T_45 == 32'h00000023;
	wire _id_ctrl_decoder_bit_T_78 = _id_ctrl_decoder_bit_T_45 == 32'h00001023;
	wire _id_ctrl_decoder_bit_T_80 = _id_ctrl_decoder_bit_T_45 == 32'h00002023;
	wire _id_ctrl_decoder_bit_T_82 = _id_ctrl_decoder_bit_T_59 == 32'h00000037;
	wire _id_ctrl_decoder_bit_T_84 = _id_ctrl_decoder_bit_T_45 == 32'h00000013;
	wire _id_ctrl_decoder_bit_T_86 = _id_ctrl_decoder_bit_T_45 == 32'h00002013;
	wire _id_ctrl_decoder_bit_T_88 = _id_ctrl_decoder_bit_T_45 == 32'h00003013;
	wire _id_ctrl_decoder_bit_T_90 = _id_ctrl_decoder_bit_T_45 == 32'h00007013;
	wire _id_ctrl_decoder_bit_T_92 = _id_ctrl_decoder_bit_T_45 == 32'h00006013;
	wire _id_ctrl_decoder_bit_T_94 = _id_ctrl_decoder_bit_T_45 == 32'h00004013;
	wire _id_ctrl_decoder_bit_T_96 = _id_ctrl_decoder_bit_T == 32'h00000033;
	wire _id_ctrl_decoder_bit_T_98 = _id_ctrl_decoder_bit_T == 32'h40000033;
	wire _id_ctrl_decoder_bit_T_100 = _id_ctrl_decoder_bit_T == 32'h00002033;
	wire _id_ctrl_decoder_bit_T_102 = _id_ctrl_decoder_bit_T == 32'h00003033;
	wire _id_ctrl_decoder_bit_T_104 = _id_ctrl_decoder_bit_T == 32'h00007033;
	wire _id_ctrl_decoder_bit_T_106 = _id_ctrl_decoder_bit_T == 32'h00006033;
	wire _id_ctrl_decoder_bit_T_108 = _id_ctrl_decoder_bit_T == 32'h00004033;
	wire _id_ctrl_decoder_bit_T_110 = _id_ctrl_decoder_bit_T == 32'h00001033;
	wire _id_ctrl_decoder_bit_T_112 = _id_ctrl_decoder_bit_T == 32'h00005033;
	wire _id_ctrl_decoder_bit_T_114 = _id_ctrl_decoder_bit_T == 32'h40005033;
	wire _id_ctrl_decoder_bit_T_116 = _id_ctrl_decoder_bit_T_45 == 32'h0000000f;
	wire _id_ctrl_decoder_bit_T_117 = ibuf_io_inst_0_bits_inst_bits == 32'h00000073;
	wire _id_ctrl_decoder_bit_T_118 = ibuf_io_inst_0_bits_inst_bits == 32'h00100073;
	wire _id_ctrl_decoder_bit_T_119 = ibuf_io_inst_0_bits_inst_bits == 32'h30200073;
	wire _id_ctrl_decoder_bit_T_120 = ibuf_io_inst_0_bits_inst_bits == 32'h10500073;
	wire _id_ctrl_decoder_bit_T_121 = ibuf_io_inst_0_bits_inst_bits == 32'h30500073;
	wire _id_ctrl_decoder_bit_T_123 = _id_ctrl_decoder_bit_T_45 == 32'h00001073;
	wire _id_ctrl_decoder_bit_T_125 = _id_ctrl_decoder_bit_T_45 == 32'h00002073;
	wire _id_ctrl_decoder_bit_T_127 = _id_ctrl_decoder_bit_T_45 == 32'h00003073;
	wire _id_ctrl_decoder_bit_T_129 = _id_ctrl_decoder_bit_T_45 == 32'h00005073;
	wire _id_ctrl_decoder_bit_T_131 = _id_ctrl_decoder_bit_T_45 == 32'h00006073;
	wire _id_ctrl_decoder_bit_T_133 = _id_ctrl_decoder_bit_T_45 == 32'h00007073;
	wire _id_ctrl_decoder_bit_T_164 = (((((((((((((((((((((((((((((_id_ctrl_decoder_bit_T_1 | _id_ctrl_decoder_bit_T_3) | _id_ctrl_decoder_bit_T_5) | _id_ctrl_decoder_bit_T_7) | _id_ctrl_decoder_bit_T_9) | _id_ctrl_decoder_bit_T_11) | _id_ctrl_decoder_bit_T_13) | _id_ctrl_decoder_bit_T_15) | _id_ctrl_decoder_bit_T_17) | _id_ctrl_decoder_bit_T_19) | _id_ctrl_decoder_bit_T_21) | _id_ctrl_decoder_bit_T_23) | _id_ctrl_decoder_bit_T_25) | _id_ctrl_decoder_bit_T_27) | _id_ctrl_decoder_bit_T_29) | _id_ctrl_decoder_bit_T_31) | _id_ctrl_decoder_bit_T_33) | _id_ctrl_decoder_bit_T_35) | _id_ctrl_decoder_bit_T_37) | _id_ctrl_decoder_bit_T_39) | _id_ctrl_decoder_bit_T_41) | _id_ctrl_decoder_bit_T_43) | _id_ctrl_decoder_bit_T_44) | _id_ctrl_decoder_bit_T_46) | _id_ctrl_decoder_bit_T_48) | _id_ctrl_decoder_bit_T_50) | _id_ctrl_decoder_bit_T_52) | _id_ctrl_decoder_bit_T_54) | _id_ctrl_decoder_bit_T_56) | _id_ctrl_decoder_bit_T_58) | _id_ctrl_decoder_bit_T_60;
	wire _id_ctrl_decoder_bit_T_194 = (((((((((((((((((((((((((((((_id_ctrl_decoder_bit_T_164 | _id_ctrl_decoder_bit_T_62) | _id_ctrl_decoder_bit_T_64) | _id_ctrl_decoder_bit_T_66) | _id_ctrl_decoder_bit_T_68) | _id_ctrl_decoder_bit_T_70) | _id_ctrl_decoder_bit_T_72) | _id_ctrl_decoder_bit_T_74) | _id_ctrl_decoder_bit_T_76) | _id_ctrl_decoder_bit_T_78) | _id_ctrl_decoder_bit_T_80) | _id_ctrl_decoder_bit_T_82) | _id_ctrl_decoder_bit_T_84) | _id_ctrl_decoder_bit_T_86) | _id_ctrl_decoder_bit_T_88) | _id_ctrl_decoder_bit_T_90) | _id_ctrl_decoder_bit_T_92) | _id_ctrl_decoder_bit_T_94) | _id_ctrl_decoder_bit_T_96) | _id_ctrl_decoder_bit_T_98) | _id_ctrl_decoder_bit_T_100) | _id_ctrl_decoder_bit_T_102) | _id_ctrl_decoder_bit_T_104) | _id_ctrl_decoder_bit_T_106) | _id_ctrl_decoder_bit_T_108) | _id_ctrl_decoder_bit_T_110) | _id_ctrl_decoder_bit_T_112) | _id_ctrl_decoder_bit_T_114) | _id_ctrl_decoder_bit_T_116) | _id_ctrl_decoder_bit_T_117) | _id_ctrl_decoder_bit_T_118;
	wire id_ctrl_decoder_0 = ((((((((_id_ctrl_decoder_bit_T_194 | _id_ctrl_decoder_bit_T_119) | _id_ctrl_decoder_bit_T_120) | _id_ctrl_decoder_bit_T_121) | _id_ctrl_decoder_bit_T_123) | _id_ctrl_decoder_bit_T_125) | _id_ctrl_decoder_bit_T_127) | _id_ctrl_decoder_bit_T_129) | _id_ctrl_decoder_bit_T_131) | _id_ctrl_decoder_bit_T_133;
	wire [31:0] _id_ctrl_decoder_T = ibuf_io_inst_0_bits_inst_bits & 32'h00000054;
	wire id_ctrl_decoder_3 = _id_ctrl_decoder_T == 32'h00000040;
	wire [31:0] _id_ctrl_decoder_T_2 = ibuf_io_inst_0_bits_inst_bits & 32'h00000048;
	wire id_ctrl_decoder_4 = _id_ctrl_decoder_T_2 == 32'h00000048;
	wire [31:0] _id_ctrl_decoder_T_4 = ibuf_io_inst_0_bits_inst_bits & 32'h0000001c;
	wire id_ctrl_decoder_5 = _id_ctrl_decoder_T_4 == 32'h00000004;
	wire [31:0] _id_ctrl_decoder_T_6 = ibuf_io_inst_0_bits_inst_bits & 32'h00000070;
	wire _id_ctrl_decoder_T_7 = _id_ctrl_decoder_T_6 == 32'h00000020;
	wire [31:0] _id_ctrl_decoder_T_8 = ibuf_io_inst_0_bits_inst_bits & 32'h00000064;
	wire _id_ctrl_decoder_T_9 = _id_ctrl_decoder_T_8 == 32'h00000020;
	wire [31:0] _id_ctrl_decoder_T_10 = ibuf_io_inst_0_bits_inst_bits & 32'h00000034;
	wire _id_ctrl_decoder_T_11 = _id_ctrl_decoder_T_10 == 32'h00000020;
	wire id_ctrl_decoder_6 = (_id_ctrl_decoder_T_7 | _id_ctrl_decoder_T_9) | _id_ctrl_decoder_T_11;
	wire [31:0] _id_ctrl_decoder_T_14 = ibuf_io_inst_0_bits_inst_bits & 32'h00004004;
	wire _id_ctrl_decoder_T_15 = _id_ctrl_decoder_T_14 == 32'h00000000;
	wire [31:0] _id_ctrl_decoder_T_16 = ibuf_io_inst_0_bits_inst_bits & 32'h00000044;
	wire _id_ctrl_decoder_T_17 = _id_ctrl_decoder_T_16 == 32'h00000000;
	wire [31:0] _id_ctrl_decoder_T_18 = ibuf_io_inst_0_bits_inst_bits & 32'h00000018;
	wire _id_ctrl_decoder_T_19 = _id_ctrl_decoder_T_18 == 32'h00000000;
	wire [31:0] _id_ctrl_decoder_T_20 = ibuf_io_inst_0_bits_inst_bits & 32'h00002050;
	wire _id_ctrl_decoder_T_21 = _id_ctrl_decoder_T_20 == 32'h00002000;
	wire id_ctrl_decoder_7 = ((_id_ctrl_decoder_T_15 | _id_ctrl_decoder_T_17) | _id_ctrl_decoder_T_19) | _id_ctrl_decoder_T_21;
	wire [31:0] _id_ctrl_decoder_T_25 = ibuf_io_inst_0_bits_inst_bits & 32'h00000058;
	wire _id_ctrl_decoder_T_26 = _id_ctrl_decoder_T_25 == 32'h00000000;
	wire [31:0] _id_ctrl_decoder_T_27 = ibuf_io_inst_0_bits_inst_bits & 32'h00000020;
	wire _id_ctrl_decoder_T_28 = _id_ctrl_decoder_T_27 == 32'h00000000;
	wire [31:0] _id_ctrl_decoder_T_29 = ibuf_io_inst_0_bits_inst_bits & 32'h0000000c;
	wire _id_ctrl_decoder_T_30 = _id_ctrl_decoder_T_29 == 32'h00000004;
	wire [31:0] _id_ctrl_decoder_T_31 = ibuf_io_inst_0_bits_inst_bits & 32'h00004050;
	wire _id_ctrl_decoder_T_32 = _id_ctrl_decoder_T_31 == 32'h00004050;
	wire _id_ctrl_decoder_T_37 = (((_id_ctrl_decoder_T_26 | _id_ctrl_decoder_T_28) | _id_ctrl_decoder_T_30) | id_ctrl_decoder_4) | _id_ctrl_decoder_T_32;
	wire _id_ctrl_decoder_T_39 = _id_ctrl_decoder_T_2 == 32'h00000000;
	wire [31:0] _id_ctrl_decoder_T_40 = ibuf_io_inst_0_bits_inst_bits & 32'h00004008;
	wire _id_ctrl_decoder_T_41 = _id_ctrl_decoder_T_40 == 32'h00004000;
	wire _id_ctrl_decoder_T_44 = (_id_ctrl_decoder_T_39 | _id_ctrl_decoder_T_19) | _id_ctrl_decoder_T_41;
	wire [1:0] id_ctrl_decoder_9 = {_id_ctrl_decoder_T_44, _id_ctrl_decoder_T_37};
	wire [31:0] _id_ctrl_decoder_T_45 = ibuf_io_inst_0_bits_inst_bits & 32'h00000050;
	wire _id_ctrl_decoder_T_46 = _id_ctrl_decoder_T_45 == 32'h00000000;
	wire _id_ctrl_decoder_T_50 = ((_id_ctrl_decoder_T_15 | _id_ctrl_decoder_T_46) | _id_ctrl_decoder_T_17) | _id_ctrl_decoder_T_19;
	wire [31:0] _id_ctrl_decoder_T_51 = ibuf_io_inst_0_bits_inst_bits & 32'h00000024;
	wire _id_ctrl_decoder_T_52 = _id_ctrl_decoder_T_51 == 32'h00000004;
	wire _id_ctrl_decoder_T_54 = _id_ctrl_decoder_T_52 | id_ctrl_decoder_4;
	wire [1:0] id_ctrl_decoder_10 = {_id_ctrl_decoder_T_54, _id_ctrl_decoder_T_50};
	wire [31:0] _id_ctrl_decoder_T_55 = ibuf_io_inst_0_bits_inst_bits & 32'h00000008;
	wire _id_ctrl_decoder_T_56 = _id_ctrl_decoder_T_55 == 32'h00000008;
	wire _id_ctrl_decoder_T_58 = _id_ctrl_decoder_T_16 == 32'h00000040;
	wire _id_ctrl_decoder_T_60 = _id_ctrl_decoder_T_56 | _id_ctrl_decoder_T_58;
	wire _id_ctrl_decoder_T_62 = _id_ctrl_decoder_T_16 == 32'h00000004;
	wire _id_ctrl_decoder_T_64 = _id_ctrl_decoder_T_62 | _id_ctrl_decoder_T_56;
	wire [31:0] _id_ctrl_decoder_T_65 = ibuf_io_inst_0_bits_inst_bits & 32'h00000014;
	wire _id_ctrl_decoder_T_66 = _id_ctrl_decoder_T_65 == 32'h00000010;
	wire [31:0] _id_ctrl_decoder_T_67 = ibuf_io_inst_0_bits_inst_bits & 32'h00000030;
	wire _id_ctrl_decoder_T_68 = _id_ctrl_decoder_T_67 == 32'h00000000;
	wire _id_ctrl_decoder_T_71 = (id_ctrl_decoder_5 | _id_ctrl_decoder_T_66) | _id_ctrl_decoder_T_68;
	wire [2:0] id_ctrl_decoder_11 = {_id_ctrl_decoder_T_71, _id_ctrl_decoder_T_64, _id_ctrl_decoder_T_60};
	wire [31:0] _id_ctrl_decoder_T_74 = ibuf_io_inst_0_bits_inst_bits & 32'h00003054;
	wire _id_ctrl_decoder_T_75 = _id_ctrl_decoder_T_74 == 32'h00001010;
	wire [31:0] _id_ctrl_decoder_T_76 = ibuf_io_inst_0_bits_inst_bits & 32'h00001058;
	wire _id_ctrl_decoder_T_77 = _id_ctrl_decoder_T_76 == 32'h00001040;
	wire [31:0] _id_ctrl_decoder_T_78 = ibuf_io_inst_0_bits_inst_bits & 32'h00007044;
	wire _id_ctrl_decoder_T_79 = _id_ctrl_decoder_T_78 == 32'h00007000;
	wire [31:0] _id_ctrl_decoder_T_80 = ibuf_io_inst_0_bits_inst_bits & 32'h02001074;
	wire _id_ctrl_decoder_T_81 = _id_ctrl_decoder_T_80 == 32'h02001030;
	wire _id_ctrl_decoder_T_85 = ((_id_ctrl_decoder_T_75 | _id_ctrl_decoder_T_77) | _id_ctrl_decoder_T_79) | _id_ctrl_decoder_T_81;
	wire [31:0] _id_ctrl_decoder_T_86 = ibuf_io_inst_0_bits_inst_bits & 32'h00004054;
	wire _id_ctrl_decoder_T_87 = _id_ctrl_decoder_T_86 == 32'h00000040;
	wire [31:0] _id_ctrl_decoder_T_88 = ibuf_io_inst_0_bits_inst_bits & 32'h00003044;
	wire _id_ctrl_decoder_T_89 = _id_ctrl_decoder_T_88 == 32'h00003000;
	wire [31:0] _id_ctrl_decoder_T_90 = ibuf_io_inst_0_bits_inst_bits & 32'h00006044;
	wire _id_ctrl_decoder_T_91 = _id_ctrl_decoder_T_90 == 32'h00006000;
	wire [31:0] _id_ctrl_decoder_T_92 = ibuf_io_inst_0_bits_inst_bits & 32'h00006018;
	wire _id_ctrl_decoder_T_93 = _id_ctrl_decoder_T_92 == 32'h00006000;
	wire [31:0] _id_ctrl_decoder_T_94 = ibuf_io_inst_0_bits_inst_bits & 32'h02002074;
	wire _id_ctrl_decoder_T_95 = _id_ctrl_decoder_T_94 == 32'h02002030;
	wire [31:0] _id_ctrl_decoder_T_96 = ibuf_io_inst_0_bits_inst_bits & 32'h40003034;
	wire _id_ctrl_decoder_T_97 = _id_ctrl_decoder_T_96 == 32'h40000030;
	wire [31:0] _id_ctrl_decoder_T_98 = ibuf_io_inst_0_bits_inst_bits & 32'h40001054;
	wire _id_ctrl_decoder_T_99 = _id_ctrl_decoder_T_98 == 32'h40001010;
	wire _id_ctrl_decoder_T_106 = (((((_id_ctrl_decoder_T_87 | _id_ctrl_decoder_T_89) | _id_ctrl_decoder_T_91) | _id_ctrl_decoder_T_93) | _id_ctrl_decoder_T_95) | _id_ctrl_decoder_T_97) | _id_ctrl_decoder_T_99;
	wire [31:0] _id_ctrl_decoder_T_107 = ibuf_io_inst_0_bits_inst_bits & 32'h02002054;
	wire _id_ctrl_decoder_T_108 = _id_ctrl_decoder_T_107 == 32'h00002010;
	wire [31:0] _id_ctrl_decoder_T_109 = ibuf_io_inst_0_bits_inst_bits & 32'h00002034;
	wire _id_ctrl_decoder_T_110 = _id_ctrl_decoder_T_109 == 32'h00002010;
	wire [31:0] _id_ctrl_decoder_T_111 = ibuf_io_inst_0_bits_inst_bits & 32'h40004054;
	wire _id_ctrl_decoder_T_112 = _id_ctrl_decoder_T_111 == 32'h00004010;
	wire [31:0] _id_ctrl_decoder_T_113 = ibuf_io_inst_0_bits_inst_bits & 32'h00005054;
	wire _id_ctrl_decoder_T_114 = _id_ctrl_decoder_T_113 == 32'h00004010;
	wire [31:0] _id_ctrl_decoder_T_115 = ibuf_io_inst_0_bits_inst_bits & 32'h00004058;
	wire _id_ctrl_decoder_T_116 = _id_ctrl_decoder_T_115 == 32'h00004040;
	wire _id_ctrl_decoder_T_121 = (((_id_ctrl_decoder_T_108 | _id_ctrl_decoder_T_110) | _id_ctrl_decoder_T_112) | _id_ctrl_decoder_T_114) | _id_ctrl_decoder_T_116;
	wire [31:0] _id_ctrl_decoder_T_122 = ibuf_io_inst_0_bits_inst_bits & 32'h02006054;
	wire _id_ctrl_decoder_T_123 = _id_ctrl_decoder_T_122 == 32'h00002010;
	wire [31:0] _id_ctrl_decoder_T_124 = ibuf_io_inst_0_bits_inst_bits & 32'h00006034;
	wire _id_ctrl_decoder_T_125 = _id_ctrl_decoder_T_124 == 32'h00002010;
	wire [31:0] _id_ctrl_decoder_T_126 = ibuf_io_inst_0_bits_inst_bits & 32'h40003054;
	wire _id_ctrl_decoder_T_127 = _id_ctrl_decoder_T_126 == 32'h40001010;
	wire _id_ctrl_decoder_T_132 = (((_id_ctrl_decoder_T_123 | _id_ctrl_decoder_T_125) | _id_ctrl_decoder_T_116) | _id_ctrl_decoder_T_97) | _id_ctrl_decoder_T_127;
	wire [3:0] id_ctrl_decoder_13 = {_id_ctrl_decoder_T_132, _id_ctrl_decoder_T_121, _id_ctrl_decoder_T_106, _id_ctrl_decoder_T_85};
	wire id_ctrl_decoder_14 = (((((((((((((((((_id_ctrl_decoder_bit_T_17 | _id_ctrl_decoder_bit_T_19) | _id_ctrl_decoder_bit_T_21) | _id_ctrl_decoder_bit_T_23) | _id_ctrl_decoder_bit_T_25) | _id_ctrl_decoder_bit_T_27) | _id_ctrl_decoder_bit_T_29) | _id_ctrl_decoder_bit_T_31) | _id_ctrl_decoder_bit_T_33) | _id_ctrl_decoder_bit_T_35) | _id_ctrl_decoder_bit_T_37) | _id_ctrl_decoder_bit_T_66) | _id_ctrl_decoder_bit_T_68) | _id_ctrl_decoder_bit_T_70) | _id_ctrl_decoder_bit_T_72) | _id_ctrl_decoder_bit_T_74) | _id_ctrl_decoder_bit_T_76) | _id_ctrl_decoder_bit_T_78) | _id_ctrl_decoder_bit_T_80;
	wire [31:0] _id_ctrl_decoder_T_133 = ibuf_io_inst_0_bits_inst_bits & 32'h00000028;
	wire _id_ctrl_decoder_T_134 = _id_ctrl_decoder_T_133 == 32'h00000020;
	wire [31:0] _id_ctrl_decoder_T_135 = ibuf_io_inst_0_bits_inst_bits & 32'h18000020;
	wire _id_ctrl_decoder_T_136 = _id_ctrl_decoder_T_135 == 32'h18000020;
	wire [31:0] _id_ctrl_decoder_T_137 = ibuf_io_inst_0_bits_inst_bits & 32'h20000020;
	wire _id_ctrl_decoder_T_138 = _id_ctrl_decoder_T_137 == 32'h20000020;
	wire _id_ctrl_decoder_T_141 = (_id_ctrl_decoder_T_134 | _id_ctrl_decoder_T_136) | _id_ctrl_decoder_T_138;
	wire [31:0] _id_ctrl_decoder_T_142 = ibuf_io_inst_0_bits_inst_bits & 32'h10000008;
	wire _id_ctrl_decoder_T_143 = _id_ctrl_decoder_T_142 == 32'h10000008;
	wire [31:0] _id_ctrl_decoder_T_144 = ibuf_io_inst_0_bits_inst_bits & 32'h40000008;
	wire _id_ctrl_decoder_T_145 = _id_ctrl_decoder_T_144 == 32'h40000008;
	wire _id_ctrl_decoder_T_147 = _id_ctrl_decoder_T_143 | _id_ctrl_decoder_T_145;
	wire [31:0] _id_ctrl_decoder_T_148 = ibuf_io_inst_0_bits_inst_bits & 32'h08000008;
	wire _id_ctrl_decoder_T_149 = _id_ctrl_decoder_T_148 == 32'h08000008;
	wire [31:0] _id_ctrl_decoder_T_150 = ibuf_io_inst_0_bits_inst_bits & 32'h80000008;
	wire _id_ctrl_decoder_T_151 = _id_ctrl_decoder_T_150 == 32'h80000008;
	wire _id_ctrl_decoder_T_154 = (_id_ctrl_decoder_T_149 | _id_ctrl_decoder_T_143) | _id_ctrl_decoder_T_151;
	wire [31:0] _id_ctrl_decoder_T_155 = ibuf_io_inst_0_bits_inst_bits & 32'h18000008;
	wire _id_ctrl_decoder_T_156 = _id_ctrl_decoder_T_155 == 32'h00000008;
	wire [4:0] id_ctrl_decoder_15 = {1'h0, _id_ctrl_decoder_T_156, _id_ctrl_decoder_T_154, _id_ctrl_decoder_T_147, _id_ctrl_decoder_T_141};
	wire [31:0] _id_ctrl_decoder_T_158 = ibuf_io_inst_0_bits_inst_bits & 32'h02000074;
	wire id_ctrl_decoder_21 = _id_ctrl_decoder_T_158 == 32'h02000030;
	wire _id_ctrl_decoder_T_161 = _id_ctrl_decoder_T_133 == 32'h00000000;
	wire _id_ctrl_decoder_T_163 = _id_ctrl_decoder_T_45 == 32'h00000010;
	wire [31:0] _id_ctrl_decoder_T_164 = ibuf_io_inst_0_bits_inst_bits & 32'h00001010;
	wire _id_ctrl_decoder_T_165 = _id_ctrl_decoder_T_164 == 32'h00001010;
	wire [31:0] _id_ctrl_decoder_T_166 = ibuf_io_inst_0_bits_inst_bits & 32'h00002008;
	wire _id_ctrl_decoder_T_167 = _id_ctrl_decoder_T_166 == 32'h00002008;
	wire [31:0] _id_ctrl_decoder_T_168 = ibuf_io_inst_0_bits_inst_bits & 32'h00002010;
	wire _id_ctrl_decoder_T_169 = _id_ctrl_decoder_T_168 == 32'h00002010;
	wire id_ctrl_decoder_22 = (((((_id_ctrl_decoder_T_161 | _id_ctrl_decoder_T_30) | _id_ctrl_decoder_T_163) | id_ctrl_decoder_4) | _id_ctrl_decoder_T_165) | _id_ctrl_decoder_T_167) | _id_ctrl_decoder_T_169;
	wire [31:0] _id_ctrl_decoder_T_176 = ibuf_io_inst_0_bits_inst_bits & 32'h00001050;
	wire _id_ctrl_decoder_T_177 = _id_ctrl_decoder_T_176 == 32'h00001050;
	wire _id_ctrl_decoder_T_180 = _id_ctrl_decoder_T_20 == 32'h00002050;
	wire _id_ctrl_decoder_T_183 = _id_ctrl_decoder_T_45 == 32'h00000050;
	wire [2:0] id_ctrl_decoder_23 = {_id_ctrl_decoder_T_183, _id_ctrl_decoder_T_180, _id_ctrl_decoder_T_177};
	wire [31:0] _id_ctrl_decoder_T_185 = ibuf_io_inst_0_bits_inst_bits & 32'h00001048;
	wire id_ctrl_decoder_24 = _id_ctrl_decoder_T_185 == 32'h00001008;
	wire [31:0] _id_ctrl_decoder_T_187 = ibuf_io_inst_0_bits_inst_bits & 32'h00002048;
	wire id_ctrl_decoder_25 = _id_ctrl_decoder_T_187 == 32'h00000008;
	wire id_ctrl_decoder_26 = _id_ctrl_decoder_T_187 == 32'h00002008;
	wire [4:0] id_raddr2 = ibuf_io_inst_0_bits_inst_rs2;
	wire [4:0] id_raddr1 = ibuf_io_inst_0_bits_inst_rs1;
	wire [4:0] id_waddr = ibuf_io_inst_0_bits_inst_rd;
	reg id_reg_fence;
	wire [31:0] _id_rs_T_4 = rf_id_rs_MPORT_data;
	wire [31:0] _id_rs_T_9 = rf_id_rs_MPORT_1_data;
	wire _id_csr_en_T = id_ctrl_decoder_23 == 3'h6;
	wire _id_csr_en_T_1 = id_ctrl_decoder_23 == 3'h7;
	wire _id_csr_en_T_2 = id_ctrl_decoder_23 == 3'h5;
	wire _id_csr_en_T_3 = _id_csr_en_T | _id_csr_en_T_1;
	wire id_csr_en = (_id_csr_en_T | _id_csr_en_T_1) | _id_csr_en_T_2;
	wire id_system_insn = id_ctrl_decoder_23 == 3'h4;
	wire id_csr_ren = _id_csr_en_T_3 & (ibuf_io_inst_0_bits_inst_rs1 == 5'h00);
	wire _id_csr_flush_T = ~id_csr_ren;
	wire id_csr_flush = id_system_insn | ((id_csr_en & ~id_csr_ren) & csr_io_decode_0_write_flush);
	wire _id_illegal_insn_T_4 = id_ctrl_decoder_21 & ~csr_io_status_isa[12];
	wire _id_illegal_insn_T_5 = ~id_ctrl_decoder_0 | _id_illegal_insn_T_4;
	wire _id_illegal_insn_T_8 = id_ctrl_decoder_26 & ~csr_io_status_isa[0];
	wire _id_illegal_insn_T_9 = _id_illegal_insn_T_5 | _id_illegal_insn_T_8;
	wire _id_illegal_insn_T_18 = ~csr_io_status_isa[2];
	wire _id_illegal_insn_T_19 = ibuf_io_inst_0_bits_rvc & ~csr_io_status_isa[2];
	wire _id_illegal_insn_T_20 = _id_illegal_insn_T_9 | _id_illegal_insn_T_19;
	wire _id_illegal_insn_T_42 = id_csr_en & (csr_io_decode_0_read_illegal | (_id_csr_flush_T & csr_io_decode_0_write_illegal));
	wire _id_illegal_insn_T_43 = _id_illegal_insn_T_20 | _id_illegal_insn_T_42;
	wire _id_illegal_insn_T_46 = ~ibuf_io_inst_0_bits_rvc & (id_system_insn & csr_io_decode_0_system_illegal);
	wire id_illegal_insn = _id_illegal_insn_T_43 | _id_illegal_insn_T_46;
	wire id_amo_aq = ibuf_io_inst_0_bits_inst_bits[26];
	wire id_amo_rl = ibuf_io_inst_0_bits_inst_bits[25];
	wire [3:0] id_fence_succ = ibuf_io_inst_0_bits_inst_bits[23:20];
	wire id_fence_next = id_ctrl_decoder_25 | (id_ctrl_decoder_26 & id_amo_aq);
	wire id_mem_busy = ~io_dmem_ordered | io_dmem_req_valid;
	wire _GEN_0 = (~id_mem_busy ? 1'h0 : id_reg_fence);
	wire id_do_fence_x9 = id_mem_busy & (((id_ctrl_decoder_26 & id_amo_rl) | id_ctrl_decoder_24) | (id_reg_fence & id_ctrl_decoder_14));
	wire id_xcpt = ((((((csr_io_interrupt | bpu_io_debug_if) | bpu_io_xcpt_if) | ibuf_io_inst_0_bits_xcpt0_ae_inst) | ibuf_io_inst_0_bits_xcpt1_pf_inst) | ibuf_io_inst_0_bits_xcpt1_gf_inst) | ibuf_io_inst_0_bits_xcpt1_ae_inst) | id_illegal_insn;
	wire [4:0] _T_11 = (ibuf_io_inst_0_bits_xcpt1_ae_inst ? 5'h01 : 5'h02);
	wire [4:0] _T_12 = (ibuf_io_inst_0_bits_xcpt1_gf_inst ? 5'h14 : _T_11);
	wire [4:0] _T_13 = (ibuf_io_inst_0_bits_xcpt1_pf_inst ? 5'h0c : _T_12);
	wire [4:0] _T_14 = (ibuf_io_inst_0_bits_xcpt0_ae_inst ? 5'h01 : _T_13);
	wire [4:0] _T_17 = (bpu_io_xcpt_if ? 5'h03 : _T_14);
	wire [4:0] _T_18 = (bpu_io_debug_if ? 5'h0e : _T_17);
	wire [4:0] ex_waddr = ex_reg_inst[11:7];
	wire [4:0] mem_waddr = mem_reg_inst[11:7];
	wire [4:0] wb_waddr = wb_reg_inst[11:7];
	wire _T_27 = ex_reg_valid & ex_ctrl_wxd;
	wire _T_28 = mem_reg_valid & mem_ctrl_wxd;
	wire _T_30 = (mem_reg_valid & mem_ctrl_wxd) & ~mem_ctrl_mem;
	wire id_bypass_src_0_0 = 5'h00 == id_raddr1;
	wire id_bypass_src_0_1 = _T_27 & (ex_waddr == id_raddr1);
	wire id_bypass_src_0_2 = _T_30 & (mem_waddr == id_raddr1);
	wire id_bypass_src_0_3 = _T_28 & (mem_waddr == id_raddr1);
	wire id_bypass_src_1_0 = 5'h00 == id_raddr2;
	wire id_bypass_src_1_1 = _T_27 & (ex_waddr == id_raddr2);
	wire id_bypass_src_1_2 = _T_30 & (mem_waddr == id_raddr2);
	wire id_bypass_src_1_3 = _T_28 & (mem_waddr == id_raddr2);
	reg ex_reg_rs_bypass_0;
	reg ex_reg_rs_bypass_1;
	reg [1:0] ex_reg_rs_lsb_0;
	reg [1:0] ex_reg_rs_lsb_1;
	reg [29:0] ex_reg_rs_msb_0;
	reg [29:0] ex_reg_rs_msb_1;
	wire [31:0] _ex_rs_T_1 = (ex_reg_rs_lsb_0 == 2'h1 ? mem_reg_wdata : 32'h00000000);
	wire [31:0] _ex_rs_T_3 = (ex_reg_rs_lsb_0 == 2'h2 ? wb_reg_wdata : _ex_rs_T_1);
	wire [31:0] _ex_rs_T_5 = (ex_reg_rs_lsb_0 == 2'h3 ? io_dmem_resp_bits_data_word_bypass : _ex_rs_T_3);
	wire [31:0] _ex_rs_T_6 = {ex_reg_rs_msb_0, ex_reg_rs_lsb_0};
	wire [31:0] _ex_rs_T_8 = (ex_reg_rs_lsb_1 == 2'h1 ? mem_reg_wdata : 32'h00000000);
	wire [31:0] _ex_rs_T_10 = (ex_reg_rs_lsb_1 == 2'h2 ? wb_reg_wdata : _ex_rs_T_8);
	wire [31:0] _ex_rs_T_12 = (ex_reg_rs_lsb_1 == 2'h3 ? io_dmem_resp_bits_data_word_bypass : _ex_rs_T_10);
	wire [31:0] _ex_rs_T_13 = {ex_reg_rs_msb_1, ex_reg_rs_lsb_1};
	wire [31:0] ex_rs_1 = (ex_reg_rs_bypass_1 ? _ex_rs_T_12 : _ex_rs_T_13);
	wire _ex_imm_sign_T = ex_ctrl_sel_imm == 3'h5;
	wire _ex_imm_sign_T_2 = ex_reg_inst[31];
	wire ex_imm_sign = (ex_ctrl_sel_imm == 3'h5 ? $signed(1'sh0) : $signed(_ex_imm_sign_T_2));
	wire _ex_imm_b30_20_T = ex_ctrl_sel_imm == 3'h2;
	wire [10:0] _ex_imm_b30_20_T_2 = ex_reg_inst[30:20];
	wire [7:0] _ex_imm_b19_12_T_4 = ex_reg_inst[19:12];
	wire _ex_imm_b11_T_2 = _ex_imm_b30_20_T | _ex_imm_sign_T;
	wire _ex_imm_b11_T_5 = ex_reg_inst[20];
	wire _ex_imm_b11_T_6 = ex_ctrl_sel_imm == 3'h1;
	wire _ex_imm_b11_T_8 = ex_reg_inst[7];
	wire _ex_imm_b11_T_9 = (ex_ctrl_sel_imm == 3'h1 ? $signed(_ex_imm_b11_T_8) : $signed(ex_imm_sign));
	wire _ex_imm_b11_T_10 = (ex_ctrl_sel_imm == 3'h3 ? $signed(_ex_imm_b11_T_5) : $signed(_ex_imm_b11_T_9));
	wire [5:0] ex_imm_b10_5 = (_ex_imm_b11_T_2 ? 6'h00 : ex_reg_inst[30:25]);
	wire _ex_imm_b4_1_T_1 = ex_ctrl_sel_imm == 3'h0;
	wire [3:0] _ex_imm_b4_1_T_8 = (_ex_imm_sign_T ? ex_reg_inst[19:16] : ex_reg_inst[24:21]);
	wire [3:0] _ex_imm_b4_1_T_9 = ((ex_ctrl_sel_imm == 3'h0) | _ex_imm_b11_T_6 ? ex_reg_inst[11:8] : _ex_imm_b4_1_T_8);
	wire [3:0] ex_imm_b4_1 = (_ex_imm_b30_20_T ? 4'h0 : _ex_imm_b4_1_T_9);
	wire _ex_imm_b0_T_6 = _ex_imm_sign_T & ex_reg_inst[15];
	wire _ex_imm_b0_T_7 = (ex_ctrl_sel_imm == 3'h4 ? ex_reg_inst[20] : _ex_imm_b0_T_6);
	wire ex_imm_b0 = (_ex_imm_b4_1_T_1 ? ex_reg_inst[7] : _ex_imm_b0_T_7);
	wire ex_imm_hi_lo_lo = (_ex_imm_b30_20_T | _ex_imm_sign_T ? $signed(1'sh0) : $signed(_ex_imm_b11_T_10));
	wire [7:0] ex_imm_hi_lo_hi = ((ex_ctrl_sel_imm != 3'h2) & (ex_ctrl_sel_imm != 3'h3) ? $signed({8 {ex_imm_sign}}) : $signed(_ex_imm_b19_12_T_4));
	wire [10:0] ex_imm_hi_hi_lo = (ex_ctrl_sel_imm == 3'h2 ? $signed(_ex_imm_b30_20_T_2) : $signed({11 {ex_imm_sign}}));
	wire ex_imm_hi_hi_hi = (ex_ctrl_sel_imm == 3'h5 ? $signed(1'sh0) : $signed(_ex_imm_sign_T_2));
	wire [31:0] ex_imm = {ex_imm_hi_hi_hi, ex_imm_hi_hi_lo, ex_imm_hi_lo_hi, ex_imm_hi_lo_lo, ex_imm_b10_5, ex_imm_b4_1, ex_imm_b0};
	wire [31:0] _ex_op1_T = (ex_reg_rs_bypass_0 ? _ex_rs_T_5 : _ex_rs_T_6);
	wire [31:0] _ex_op1_T_3 = (2'h1 == ex_ctrl_sel_alu1 ? $signed(_ex_op1_T) : $signed(32'sh00000000));
	wire [31:0] _ex_op2_T = (ex_reg_rs_bypass_1 ? _ex_rs_T_12 : _ex_rs_T_13);
	wire [3:0] _ex_op2_T_1 = (ex_reg_rvc ? $signed(4'sh2) : $signed(4'sh4));
	wire [31:0] _ex_op2_T_3 = (2'h2 == ex_ctrl_sel_alu2 ? $signed(_ex_op2_T) : $signed(32'sh00000000));
	wire [31:0] _ex_op2_T_5 = (2'h3 == ex_ctrl_sel_alu2 ? $signed(ex_imm) : $signed(_ex_op2_T_3));
	wire _T_134 = id_raddr1 != 5'h00;
	wire _T_135 = id_ctrl_decoder_7 & (id_raddr1 != 5'h00);
	wire _data_hazard_ex_T = id_raddr1 == ex_waddr;
	wire _T_136 = id_raddr2 != 5'h00;
	wire _T_137 = id_ctrl_decoder_6 & (id_raddr2 != 5'h00);
	wire _data_hazard_ex_T_2 = id_raddr2 == ex_waddr;
	wire _T_139 = id_ctrl_decoder_22 & (id_waddr != 5'h00);
	wire _data_hazard_ex_T_4 = id_waddr == ex_waddr;
	wire _data_hazard_ex_T_7 = ((_T_135 & _data_hazard_ex_T) | (_T_137 & _data_hazard_ex_T_2)) | (_T_139 & _data_hazard_ex_T_4);
	wire data_hazard_ex = ex_ctrl_wxd & _data_hazard_ex_T_7;
	wire ex_cannot_bypass = (((ex_ctrl_csr != 3'h0) | ex_ctrl_jalr) | ex_ctrl_mem) | ex_ctrl_div;
	wire id_ex_hazard = ex_reg_valid & (data_hazard_ex & ex_cannot_bypass);
	wire _data_hazard_mem_T = id_raddr1 == mem_waddr;
	wire _data_hazard_mem_T_2 = id_raddr2 == mem_waddr;
	wire _data_hazard_mem_T_4 = id_waddr == mem_waddr;
	wire _data_hazard_mem_T_7 = ((_T_135 & _data_hazard_mem_T) | (_T_137 & _data_hazard_mem_T_2)) | (_T_139 & _data_hazard_mem_T_4);
	wire data_hazard_mem = mem_ctrl_wxd & _data_hazard_mem_T_7;
	wire mem_cannot_bypass = ((mem_ctrl_csr != 3'h0) | (mem_ctrl_mem & mem_reg_slow_bypass)) | mem_ctrl_div;
	wire id_mem_hazard = mem_reg_valid & (data_hazard_mem & mem_cannot_bypass);
	wire _data_hazard_wb_T = id_raddr1 == wb_waddr;
	wire _data_hazard_wb_T_2 = id_raddr2 == wb_waddr;
	wire _data_hazard_wb_T_4 = id_waddr == wb_waddr;
	wire _data_hazard_wb_T_7 = ((_T_135 & _data_hazard_wb_T) | (_T_137 & _data_hazard_wb_T_2)) | (_T_139 & _data_hazard_wb_T_4);
	wire data_hazard_wb = wb_ctrl_wxd & _data_hazard_wb_T_7;
	wire wb_dcache_miss = wb_ctrl_mem & ~io_dmem_resp_valid;
	wire wb_set_sboard = wb_ctrl_div | wb_dcache_miss;
	wire id_wb_hazard = wb_reg_valid & (data_hazard_wb & wb_set_sboard);
	reg [31:0] _r;
	wire [31:0] r = {_r[31:1], 1'h0};
	wire [31:0] _id_sboard_hazard_T = r >> id_raddr1;
	wire dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
	wire dmem_resp_replay = dmem_resp_valid & io_dmem_resp_bits_replay;
	wire dmem_resp_xpu = ~io_dmem_resp_bits_tag[0];
	wire ll_wen_x2 = div_io_resp_ready & div_io_resp_valid;
	wire ll_wen = (dmem_resp_replay & dmem_resp_xpu) | ll_wen_x2;
	wire [4:0] dmem_resp_waddr = io_dmem_resp_bits_tag[5:1];
	wire [4:0] ll_waddr = (dmem_resp_replay & dmem_resp_xpu ? dmem_resp_waddr : div_io_resp_bits_tag);
	wire _id_sboard_hazard_T_3 = ll_wen & (ll_waddr == id_raddr1);
	wire _id_sboard_hazard_T_5 = _id_sboard_hazard_T[0] & ~_id_sboard_hazard_T_3;
	wire [31:0] _id_sboard_hazard_T_7 = r >> id_raddr2;
	wire _id_sboard_hazard_T_10 = ll_wen & (ll_waddr == id_raddr2);
	wire _id_sboard_hazard_T_12 = _id_sboard_hazard_T_7[0] & ~_id_sboard_hazard_T_10;
	wire [31:0] _id_sboard_hazard_T_14 = r >> id_waddr;
	wire _id_sboard_hazard_T_17 = ll_wen & (ll_waddr == id_waddr);
	wire _id_sboard_hazard_T_19 = _id_sboard_hazard_T_14[0] & ~_id_sboard_hazard_T_17;
	wire id_sboard_hazard = ((_T_135 & _id_sboard_hazard_T_5) | (_T_137 & _id_sboard_hazard_T_12)) | (_T_139 & _id_sboard_hazard_T_19);
	wire _ctrl_stalld_T_5 = csr_io_singleStep & ((ex_reg_valid | mem_reg_valid) | wb_reg_valid);
	wire _ctrl_stalld_T_6 = (((id_ex_hazard | id_mem_hazard) | id_wb_hazard) | id_sboard_hazard) | _ctrl_stalld_T_5;
	reg blocked;
	wire _dcache_blocked_T = ~io_dmem_perf_grant;
	wire dcache_blocked = blocked & ~io_dmem_perf_grant;
	wire _ctrl_stalld_T_13 = id_ctrl_decoder_14 & dcache_blocked;
	wire _ctrl_stalld_T_14 = _ctrl_stalld_T_6 | _ctrl_stalld_T_13;
	wire wb_wxd = wb_reg_valid & wb_ctrl_wxd;
	wire _ctrl_stalld_T_17 = ~wb_wxd;
	wire _ctrl_stalld_T_22 = id_ctrl_decoder_21 & (~(div_io_req_ready | (div_io_resp_valid & ~wb_wxd)) | div_io_req_valid);
	wire _ctrl_stalld_T_23 = _ctrl_stalld_T_14 | _ctrl_stalld_T_22;
	wire _ctrl_stalld_T_26 = _ctrl_stalld_T_23 | id_do_fence_x9;
	wire _ctrl_stalld_T_27 = _ctrl_stalld_T_26 | csr_io_csr_stall;
	wire ctrl_stalld = _ctrl_stalld_T_27 | id_reg_pause;
	wire ctrl_killd = (((~ibuf_io_inst_0_valid | ibuf_io_inst_0_bits_replay) | take_pc_mem_wb) | ctrl_stalld) | csr_io_interrupt;
	wire _ex_reg_valid_T = ~ctrl_killd;
	wire _ex_reg_replay_T = ~take_pc_mem_wb;
	wire _ex_reg_replay_T_1 = ~take_pc_mem_wb & ibuf_io_inst_0_valid;
	wire _GEN_1 = (id_ctrl_decoder_25 & (id_fence_succ == 4'h0)) | id_reg_pause;
	wire _GEN_2 = id_fence_next | _GEN_0;
	wire [2:0] _T_35 = {ibuf_io_inst_0_bits_xcpt1_pf_inst, ibuf_io_inst_0_bits_xcpt1_gf_inst, ibuf_io_inst_0_bits_xcpt1_ae_inst};
	wire _GEN_5 = |_T_35 | ibuf_io_inst_0_bits_rvc;
	wire [2:0] _T_37 = {2'h0, ibuf_io_inst_0_bits_xcpt0_ae_inst};
	wire _T_40 = id_ctrl_decoder_15 == 5'h14;
	wire _T_41 = id_ctrl_decoder_15 == 5'h15;
	wire _T_42 = id_ctrl_decoder_15 == 5'h16;
	wire _T_43 = id_ctrl_decoder_15 == 5'h05;
	wire _T_46 = ((_T_40 | _T_41) | _T_42) | _T_43;
	wire [1:0] _ex_reg_mem_size_T_6 = {_T_136, _T_134};
	wire do_bypass = ((id_bypass_src_0_0 | id_bypass_src_0_1) | id_bypass_src_0_2) | id_bypass_src_0_3;
	wire [1:0] _bypass_src_T = (id_bypass_src_0_2 ? 2'h2 : 2'h3);
	wire [1:0] _bypass_src_T_1 = (id_bypass_src_0_1 ? 2'h1 : _bypass_src_T);
	wire wb_valid = (wb_reg_valid & ~replay_wb_common) & ~wb_xcpt;
	wire wb_wen = wb_valid & wb_ctrl_wxd;
	wire rf_wen = wb_wen | ll_wen;
	wire [4:0] rf_waddr = (ll_wen ? ll_waddr : wb_waddr);
	wire _T_129 = rf_waddr != 5'h00;
	wire _rf_wdata_T = dmem_resp_valid & dmem_resp_xpu;
	wire [31:0] ll_wdata = div_io_resp_bits_data;
	wire [31:0] _rf_wdata_T_4 = (wb_ctrl_csr != 3'h0 ? csr_io_rw_rdata : wb_reg_wdata);
	wire [31:0] _rf_wdata_T_5 = (ll_wen ? ll_wdata : _rf_wdata_T_4);
	wire [31:0] rf_wdata = (dmem_resp_valid & dmem_resp_xpu ? io_dmem_resp_bits_data : _rf_wdata_T_5);
	wire [31:0] _GEN_233 = (rf_waddr == id_raddr1 ? rf_wdata : _id_rs_T_4);
	wire [31:0] _GEN_240 = (rf_waddr != 5'h00 ? _GEN_233 : _id_rs_T_4);
	wire [31:0] id_rs_0 = (rf_wen ? _GEN_240 : _id_rs_T_4);
	wire do_bypass_1 = ((id_bypass_src_1_0 | id_bypass_src_1_1) | id_bypass_src_1_2) | id_bypass_src_1_3;
	wire [1:0] _bypass_src_T_2 = (id_bypass_src_1_2 ? 2'h2 : 2'h3);
	wire [31:0] _GEN_234 = (rf_waddr == id_raddr2 ? rf_wdata : _id_rs_T_9);
	wire [31:0] _GEN_241 = (rf_waddr != 5'h00 ? _GEN_234 : _id_rs_T_9);
	wire [31:0] id_rs_1 = (rf_wen ? _GEN_241 : _id_rs_T_9);
	wire [31:0] inst = (ibuf_io_inst_0_bits_rvc ? {16'd0, ibuf_io_inst_0_bits_raw[15:0]} : ibuf_io_inst_0_bits_raw);
	wire id_load_use = (mem_reg_valid & data_hazard_mem) & mem_ctrl_mem;
	wire ex_pc_valid = (ex_reg_valid | ex_reg_replay) | ex_reg_xcpt_interrupt;
	wire _replay_ex_structural_T = ~io_dmem_req_ready;
	wire _replay_ex_structural_T_3 = ex_ctrl_div & ~div_io_req_ready;
	wire replay_ex_structural = (ex_ctrl_mem & ~io_dmem_req_ready) | _replay_ex_structural_T_3;
	wire replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
	wire replay_ex = ex_reg_replay | (ex_reg_valid & (replay_ex_structural | replay_ex_load_use));
	wire ctrl_killx = (take_pc_mem_wb | replay_ex) | ~ex_reg_valid;
	wire _ex_slow_bypass_T = ex_ctrl_mem_cmd == 5'h07;
	wire ex_slow_bypass = (ex_ctrl_mem_cmd == 5'h07) | (ex_reg_mem_size < 2'h2);
	wire ex_xcpt = ex_reg_xcpt_interrupt | ex_reg_xcpt;
	wire mem_pc_valid = (mem_reg_valid | mem_reg_replay) | mem_reg_xcpt_interrupt;
	wire mem_br_target_sign = mem_reg_inst[31];
	wire [5:0] mem_br_target_b10_5 = mem_reg_inst[30:25];
	wire [3:0] mem_br_target_b4_1 = mem_reg_inst[11:8];
	wire mem_br_target_hi_lo_lo = mem_reg_inst[7];
	wire [7:0] mem_br_target_hi_lo_hi = {8 {mem_br_target_sign}};
	wire [10:0] mem_br_target_hi_hi_lo = {11 {mem_br_target_sign}};
	wire mem_br_target_hi_hi_hi = mem_reg_inst[31];
	wire [31:0] _mem_br_target_T_3 = {mem_br_target_hi_hi_hi, mem_br_target_hi_hi_lo, mem_br_target_hi_lo_hi, mem_br_target_hi_lo_lo, mem_br_target_b10_5, mem_br_target_b4_1, 1'h0};
	wire mem_br_target_hi_lo_lo_1 = mem_reg_inst[20];
	wire [7:0] mem_br_target_hi_lo_hi_1 = mem_reg_inst[19:12];
	wire [31:0] _mem_br_target_T_5 = {mem_br_target_hi_hi_hi, mem_br_target_hi_hi_lo, mem_br_target_hi_lo_hi_1, mem_br_target_hi_lo_lo_1, mem_br_target_b10_5, mem_reg_inst[24:21], 1'h0};
	wire [3:0] _mem_br_target_T_6 = (mem_reg_rvc ? $signed(4'sh2) : $signed(4'sh4));
	wire [31:0] _mem_br_target_T_7 = (mem_ctrl_jal ? $signed(_mem_br_target_T_5) : $signed({{28 {_mem_br_target_T_6[3]}}, _mem_br_target_T_6}));
	wire [31:0] _mem_br_target_T_8 = (_mem_cfi_taken_T ? $signed(_mem_br_target_T_3) : $signed(_mem_br_target_T_7));
	wire [31:0] mem_br_target = $signed(mem_reg_pc) + $signed(_mem_br_target_T_8);
	wire [31:0] _mem_npc_T_2 = (mem_ctrl_jalr ? $signed(mem_reg_wdata) : $signed(mem_br_target));
	wire [31:0] mem_npc = $signed(_mem_npc_T_2) & -32'sh00000002;
	wire _mem_wrong_npc_T_3 = (ibuf_io_inst_0_valid | ibuf_io_imem_valid ? mem_npc != ibuf_io_pc : 1'h1);
	wire mem_wrong_npc = (ex_pc_valid ? mem_npc != ex_reg_pc : _mem_wrong_npc_T_3);
	wire mem_npc_misaligned = _id_illegal_insn_T_18 & mem_npc[1];
	wire [31:0] mem_int_wdata = (_take_pc_mem_T & (mem_ctrl_jalr ^ mem_npc_misaligned) ? $signed(mem_br_target) : $signed(mem_reg_wdata));
	wire mem_cfi = (mem_ctrl_branch | mem_ctrl_jalr) | mem_ctrl_jal;
	wire _mem_reg_valid_T = ~ctrl_killx;
	wire _mem_reg_load_T = ex_ctrl_mem_cmd == 5'h00;
	wire _mem_reg_load_T_1 = ex_ctrl_mem_cmd == 5'h10;
	wire _mem_reg_load_T_2 = ex_ctrl_mem_cmd == 5'h06;
	wire _mem_reg_load_T_6 = ((_mem_reg_load_T | _mem_reg_load_T_1) | _mem_reg_load_T_2) | _ex_slow_bypass_T;
	wire _mem_reg_load_T_7 = ex_ctrl_mem_cmd == 5'h04;
	wire _mem_reg_load_T_8 = ex_ctrl_mem_cmd == 5'h09;
	wire _mem_reg_load_T_9 = ex_ctrl_mem_cmd == 5'h0a;
	wire _mem_reg_load_T_10 = ex_ctrl_mem_cmd == 5'h0b;
	wire _mem_reg_load_T_13 = ((_mem_reg_load_T_7 | _mem_reg_load_T_8) | _mem_reg_load_T_9) | _mem_reg_load_T_10;
	wire _mem_reg_load_T_14 = ex_ctrl_mem_cmd == 5'h08;
	wire _mem_reg_load_T_15 = ex_ctrl_mem_cmd == 5'h0c;
	wire _mem_reg_load_T_16 = ex_ctrl_mem_cmd == 5'h0d;
	wire _mem_reg_load_T_17 = ex_ctrl_mem_cmd == 5'h0e;
	wire _mem_reg_load_T_18 = ex_ctrl_mem_cmd == 5'h0f;
	wire _mem_reg_load_T_22 = (((_mem_reg_load_T_14 | _mem_reg_load_T_15) | _mem_reg_load_T_16) | _mem_reg_load_T_17) | _mem_reg_load_T_18;
	wire _mem_reg_load_T_23 = _mem_reg_load_T_13 | _mem_reg_load_T_22;
	wire _mem_reg_load_T_24 = _mem_reg_load_T_6 | _mem_reg_load_T_23;
	wire _mem_reg_store_T_22 = (((ex_ctrl_mem_cmd == 5'h01) | (ex_ctrl_mem_cmd == 5'h11)) | _ex_slow_bypass_T) | _mem_reg_load_T_23;
	wire [31:0] _mem_reg_wdata_T = alu_io_out;
	wire [31:0] _mem_reg_rs2_T_3 = {ex_rs_1[7:0], ex_rs_1[7:0], ex_rs_1[7:0], ex_rs_1[7:0]};
	wire [31:0] _mem_reg_rs2_T_6 = {ex_rs_1[15:0], ex_rs_1[15:0]};
	wire [31:0] _mem_reg_rs2_T_7 = (ex_reg_mem_size == 2'h1 ? _mem_reg_rs2_T_6 : ex_rs_1);
	wire _GEN_79 = (ex_ctrl_jalr & csr_io_status_debug) | ex_ctrl_fence_i;
	wire _GEN_80 = (ex_ctrl_jalr & csr_io_status_debug) | ex_reg_flush_pipe;
	wire mem_breakpoint = (mem_reg_load & bpu_io_xcpt_ld) | (mem_reg_store & bpu_io_xcpt_st);
	wire mem_debug_breakpoint = (mem_reg_load & bpu_io_debug_ld) | (mem_reg_store & bpu_io_debug_st);
	wire mem_ldst_xcpt = mem_debug_breakpoint | mem_breakpoint;
	wire [3:0] mem_ldst_cause = (mem_debug_breakpoint ? 4'he : 4'h3);
	wire _T_70 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
	wire _T_71 = mem_reg_valid & mem_npc_misaligned;
	wire _T_72 = mem_reg_valid & mem_ldst_xcpt;
	wire mem_xcpt = (_T_70 | _T_71) | _T_72;
	wire [3:0] _T_74 = (_T_71 ? 4'h0 : mem_ldst_cause);
	wire dcache_kill_mem = _T_28 & io_dmem_replay_next;
	wire replay_mem = dcache_kill_mem | mem_reg_replay;
	wire killm_common = ((dcache_kill_mem | take_pc_wb) | mem_reg_xcpt) | ~mem_reg_valid;
	reg div_io_kill_REG;
	wire ctrl_killm = killm_common | mem_xcpt;
	wire _wb_reg_valid_T = ~ctrl_killm;
	wire _wb_reg_replay_T = ~take_pc_wb;
	wire [2:0] _T_113 = (_T_103 ? 3'h6 : 3'h4);
	wire [2:0] _T_114 = (_T_101 ? 3'h5 : _T_113);
	wire [2:0] _T_115 = (_T_99 ? 3'h7 : _T_114);
	wire [4:0] _T_116 = {2'd0, _T_115};
	wire [4:0] _T_118 = (_T_93 ? 5'h0d : _T_116);
	wire [4:0] _T_119 = (_T_91 ? 5'h0f : _T_118);
	wire [15:0] _csr_io_inst_0_T_3 = (&wb_reg_raw_inst[1:0] ? wb_reg_inst[31:16] : 16'h0000);
	wire [31:0] _io_fpu_time_T = csr_io_time;
	wire tval_dmem_addr = ~wb_reg_xcpt;
	wire _tval_any_addr_T = wb_reg_cause == 32'h00000003;
	wire _tval_any_addr_T_1 = wb_reg_cause == 32'h00000001;
	wire _tval_any_addr_T_2 = wb_reg_cause == 32'h0000000c;
	wire _tval_any_addr_T_3 = wb_reg_cause == 32'h00000014;
	wire _tval_any_addr_T_6 = ((_tval_any_addr_T | _tval_any_addr_T_1) | _tval_any_addr_T_2) | _tval_any_addr_T_3;
	wire tval_any_addr = tval_dmem_addr | _tval_any_addr_T_6;
	wire tval_inst = wb_reg_cause == 32'h00000002;
	wire tval_valid = wb_xcpt & (tval_any_addr | tval_inst);
	wire htval_valid_imem = wb_reg_xcpt & _tval_any_addr_T_3;
	wire _csr_io_htval_T_3 = ~reset;
	wire [2:0] _csr_io_rw_cmd_T = (wb_reg_valid ? 3'h0 : 3'h4);
	wire [2:0] _csr_io_rw_cmd_T_1 = ~_csr_io_rw_cmd_T;
	wire [31:0] _T_140 = 32'h00000001 << ll_waddr;
	wire [31:0] _T_141 = (ll_wen ? _T_140 : 32'h00000000);
	wire [31:0] _T_142 = ~_T_141;
	wire [31:0] _T_143 = r & _T_142;
	wire _T_145 = wb_set_sboard & wb_wen;
	wire [31:0] _T_146 = 32'h00000001 << wb_waddr;
	wire [31:0] _T_147 = (_T_145 ? _T_146 : 32'h00000000);
	wire [31:0] _T_148 = _T_143 | _T_147;
	wire _T_149 = ll_wen | _T_145;
	wire [31:0] _io_imem_req_bits_pc_T_1 = (replay_wb_common ? wb_reg_pc : mem_npc);
	wire [5:0] ex_dcache_tag = {ex_waddr, 1'h0};
	wire unpause = ((csr_io_time[4:0] == 5'h00) | csr_io_inhibit_cycle) | take_pc_mem_wb;
	wire coreMonitorBundle_valid = csr_io_trace_0_valid & ~csr_io_trace_0_exception;
	wire [31:0] coreMonitorBundle_pc = csr_io_trace_0_iaddr;
	wire coreMonitorBundle_wrenx = wb_wen & ~wb_set_sboard;
	reg [31:0] coreMonitorBundle_rd0val_x23;
	reg [31:0] coreMonitorBundle_rd0val_REG;
	reg [31:0] coreMonitorBundle_rd1val_x29;
	reg [31:0] coreMonitorBundle_rd1val_REG;
	wire [4:0] _T_151 = (wb_ctrl_wxd ? wb_waddr : 5'h00);
	wire [31:0] _T_152 = (coreMonitorBundle_wrenx ? rf_wdata : 32'h00000000);
	wire [4:0] _T_154 = (wb_ctrl_rxs1 ? wb_reg_inst[19:15] : 5'h00);
	wire [31:0] _T_156 = (wb_ctrl_rxs1 ? coreMonitorBundle_rd0val_REG : 32'h00000000);
	wire [4:0] _T_158 = (wb_ctrl_rxs2 ? wb_reg_inst[24:20] : 5'h00);
	wire [31:0] _T_160 = (wb_ctrl_rxs2 ? coreMonitorBundle_rd1val_REG : 32'h00000000);
	wire [31:0] coreMonitorBundle_inst = csr_io_trace_0_insn;
	IBuf ibuf(
		.clock(ibuf_clock),
		.reset(ibuf_reset),
		.io_imem_ready(ibuf_io_imem_ready),
		.io_imem_valid(ibuf_io_imem_valid),
		.io_imem_bits_pc(ibuf_io_imem_bits_pc),
		.io_imem_bits_data(ibuf_io_imem_bits_data),
		.io_imem_bits_xcpt_ae_inst(ibuf_io_imem_bits_xcpt_ae_inst),
		.io_imem_bits_replay(ibuf_io_imem_bits_replay),
		.io_kill(ibuf_io_kill),
		.io_pc(ibuf_io_pc),
		.io_inst_0_ready(ibuf_io_inst_0_ready),
		.io_inst_0_valid(ibuf_io_inst_0_valid),
		.io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),
		.io_inst_0_bits_xcpt1_pf_inst(ibuf_io_inst_0_bits_xcpt1_pf_inst),
		.io_inst_0_bits_xcpt1_gf_inst(ibuf_io_inst_0_bits_xcpt1_gf_inst),
		.io_inst_0_bits_xcpt1_ae_inst(ibuf_io_inst_0_bits_xcpt1_ae_inst),
		.io_inst_0_bits_replay(ibuf_io_inst_0_bits_replay),
		.io_inst_0_bits_rvc(ibuf_io_inst_0_bits_rvc),
		.io_inst_0_bits_inst_bits(ibuf_io_inst_0_bits_inst_bits),
		.io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
		.io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
		.io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
		.io_inst_0_bits_raw(ibuf_io_inst_0_bits_raw)
	);
	CSRFile csr(
		.clock(csr_clock),
		.reset(csr_reset),
		.io_ungated_clock(csr_io_ungated_clock),
		.io_interrupts_debug(csr_io_interrupts_debug),
		.io_interrupts_mtip(csr_io_interrupts_mtip),
		.io_interrupts_msip(csr_io_interrupts_msip),
		.io_interrupts_meip(csr_io_interrupts_meip),
		.io_hartid(csr_io_hartid),
		.io_rw_addr(csr_io_rw_addr),
		.io_rw_cmd(csr_io_rw_cmd),
		.io_rw_rdata(csr_io_rw_rdata),
		.io_rw_wdata(csr_io_rw_wdata),
		.io_decode_0_inst(csr_io_decode_0_inst),
		.io_decode_0_fp_illegal(csr_io_decode_0_fp_illegal),
		.io_decode_0_fp_csr(csr_io_decode_0_fp_csr),
		.io_decode_0_read_illegal(csr_io_decode_0_read_illegal),
		.io_decode_0_write_illegal(csr_io_decode_0_write_illegal),
		.io_decode_0_write_flush(csr_io_decode_0_write_flush),
		.io_decode_0_system_illegal(csr_io_decode_0_system_illegal),
		.io_csr_stall(csr_io_csr_stall),
		.io_eret(csr_io_eret),
		.io_singleStep(csr_io_singleStep),
		.io_status_debug(csr_io_status_debug),
		.io_status_cease(csr_io_status_cease),
		.io_status_wfi(csr_io_status_wfi),
		.io_status_isa(csr_io_status_isa),
		.io_status_dprv(csr_io_status_dprv),
		.io_status_dv(csr_io_status_dv),
		.io_status_prv(csr_io_status_prv),
		.io_status_v(csr_io_status_v),
		.io_status_sd(csr_io_status_sd),
		.io_status_zero2(csr_io_status_zero2),
		.io_status_mpv(csr_io_status_mpv),
		.io_status_gva(csr_io_status_gva),
		.io_status_mbe(csr_io_status_mbe),
		.io_status_sbe(csr_io_status_sbe),
		.io_status_sxl(csr_io_status_sxl),
		.io_status_uxl(csr_io_status_uxl),
		.io_status_sd_rv32(csr_io_status_sd_rv32),
		.io_status_zero1(csr_io_status_zero1),
		.io_status_tsr(csr_io_status_tsr),
		.io_status_tw(csr_io_status_tw),
		.io_status_tvm(csr_io_status_tvm),
		.io_status_mxr(csr_io_status_mxr),
		.io_status_sum(csr_io_status_sum),
		.io_status_mprv(csr_io_status_mprv),
		.io_status_xs(csr_io_status_xs),
		.io_status_fs(csr_io_status_fs),
		.io_status_mpp(csr_io_status_mpp),
		.io_status_vs(csr_io_status_vs),
		.io_status_spp(csr_io_status_spp),
		.io_status_mpie(csr_io_status_mpie),
		.io_status_ube(csr_io_status_ube),
		.io_status_spie(csr_io_status_spie),
		.io_status_upie(csr_io_status_upie),
		.io_status_mie(csr_io_status_mie),
		.io_status_hie(csr_io_status_hie),
		.io_status_sie(csr_io_status_sie),
		.io_status_uie(csr_io_status_uie),
		.io_evec(csr_io_evec),
		.io_exception(csr_io_exception),
		.io_retire(csr_io_retire),
		.io_cause(csr_io_cause),
		.io_pc(csr_io_pc),
		.io_tval(csr_io_tval),
		.io_gva(csr_io_gva),
		.io_time(csr_io_time),
		.io_interrupt(csr_io_interrupt),
		.io_interrupt_cause(csr_io_interrupt_cause),
		.io_bp_0_control_action(csr_io_bp_0_control_action),
		.io_bp_0_control_tmatch(csr_io_bp_0_control_tmatch),
		.io_bp_0_control_x(csr_io_bp_0_control_x),
		.io_bp_0_control_w(csr_io_bp_0_control_w),
		.io_bp_0_control_r(csr_io_bp_0_control_r),
		.io_bp_0_address(csr_io_bp_0_address),
		.io_pmp_0_cfg_l(csr_io_pmp_0_cfg_l),
		.io_pmp_0_cfg_a(csr_io_pmp_0_cfg_a),
		.io_pmp_0_cfg_x(csr_io_pmp_0_cfg_x),
		.io_pmp_0_cfg_w(csr_io_pmp_0_cfg_w),
		.io_pmp_0_cfg_r(csr_io_pmp_0_cfg_r),
		.io_pmp_0_addr(csr_io_pmp_0_addr),
		.io_pmp_0_mask(csr_io_pmp_0_mask),
		.io_pmp_1_cfg_l(csr_io_pmp_1_cfg_l),
		.io_pmp_1_cfg_a(csr_io_pmp_1_cfg_a),
		.io_pmp_1_cfg_x(csr_io_pmp_1_cfg_x),
		.io_pmp_1_cfg_w(csr_io_pmp_1_cfg_w),
		.io_pmp_1_cfg_r(csr_io_pmp_1_cfg_r),
		.io_pmp_1_addr(csr_io_pmp_1_addr),
		.io_pmp_1_mask(csr_io_pmp_1_mask),
		.io_pmp_2_cfg_l(csr_io_pmp_2_cfg_l),
		.io_pmp_2_cfg_a(csr_io_pmp_2_cfg_a),
		.io_pmp_2_cfg_x(csr_io_pmp_2_cfg_x),
		.io_pmp_2_cfg_w(csr_io_pmp_2_cfg_w),
		.io_pmp_2_cfg_r(csr_io_pmp_2_cfg_r),
		.io_pmp_2_addr(csr_io_pmp_2_addr),
		.io_pmp_2_mask(csr_io_pmp_2_mask),
		.io_pmp_3_cfg_l(csr_io_pmp_3_cfg_l),
		.io_pmp_3_cfg_a(csr_io_pmp_3_cfg_a),
		.io_pmp_3_cfg_x(csr_io_pmp_3_cfg_x),
		.io_pmp_3_cfg_w(csr_io_pmp_3_cfg_w),
		.io_pmp_3_cfg_r(csr_io_pmp_3_cfg_r),
		.io_pmp_3_addr(csr_io_pmp_3_addr),
		.io_pmp_3_mask(csr_io_pmp_3_mask),
		.io_pmp_4_cfg_l(csr_io_pmp_4_cfg_l),
		.io_pmp_4_cfg_a(csr_io_pmp_4_cfg_a),
		.io_pmp_4_cfg_x(csr_io_pmp_4_cfg_x),
		.io_pmp_4_cfg_w(csr_io_pmp_4_cfg_w),
		.io_pmp_4_cfg_r(csr_io_pmp_4_cfg_r),
		.io_pmp_4_addr(csr_io_pmp_4_addr),
		.io_pmp_4_mask(csr_io_pmp_4_mask),
		.io_pmp_5_cfg_l(csr_io_pmp_5_cfg_l),
		.io_pmp_5_cfg_a(csr_io_pmp_5_cfg_a),
		.io_pmp_5_cfg_x(csr_io_pmp_5_cfg_x),
		.io_pmp_5_cfg_w(csr_io_pmp_5_cfg_w),
		.io_pmp_5_cfg_r(csr_io_pmp_5_cfg_r),
		.io_pmp_5_addr(csr_io_pmp_5_addr),
		.io_pmp_5_mask(csr_io_pmp_5_mask),
		.io_pmp_6_cfg_l(csr_io_pmp_6_cfg_l),
		.io_pmp_6_cfg_a(csr_io_pmp_6_cfg_a),
		.io_pmp_6_cfg_x(csr_io_pmp_6_cfg_x),
		.io_pmp_6_cfg_w(csr_io_pmp_6_cfg_w),
		.io_pmp_6_cfg_r(csr_io_pmp_6_cfg_r),
		.io_pmp_6_addr(csr_io_pmp_6_addr),
		.io_pmp_6_mask(csr_io_pmp_6_mask),
		.io_pmp_7_cfg_l(csr_io_pmp_7_cfg_l),
		.io_pmp_7_cfg_a(csr_io_pmp_7_cfg_a),
		.io_pmp_7_cfg_x(csr_io_pmp_7_cfg_x),
		.io_pmp_7_cfg_w(csr_io_pmp_7_cfg_w),
		.io_pmp_7_cfg_r(csr_io_pmp_7_cfg_r),
		.io_pmp_7_addr(csr_io_pmp_7_addr),
		.io_pmp_7_mask(csr_io_pmp_7_mask),
		.io_inhibit_cycle(csr_io_inhibit_cycle),
		.io_inst_0(csr_io_inst_0),
		.io_trace_0_valid(csr_io_trace_0_valid),
		.io_trace_0_iaddr(csr_io_trace_0_iaddr),
		.io_trace_0_insn(csr_io_trace_0_insn),
		.io_trace_0_exception(csr_io_trace_0_exception),
		.io_customCSRs_0_value(csr_io_customCSRs_0_value)
	);
	BreakpointUnit bpu(
		.io_status_debug(bpu_io_status_debug),
		.io_bp_0_control_action(bpu_io_bp_0_control_action),
		.io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),
		.io_bp_0_control_x(bpu_io_bp_0_control_x),
		.io_bp_0_control_w(bpu_io_bp_0_control_w),
		.io_bp_0_control_r(bpu_io_bp_0_control_r),
		.io_bp_0_address(bpu_io_bp_0_address),
		.io_pc(bpu_io_pc),
		.io_ea(bpu_io_ea),
		.io_xcpt_if(bpu_io_xcpt_if),
		.io_xcpt_ld(bpu_io_xcpt_ld),
		.io_xcpt_st(bpu_io_xcpt_st),
		.io_debug_if(bpu_io_debug_if),
		.io_debug_ld(bpu_io_debug_ld),
		.io_debug_st(bpu_io_debug_st)
	);
	ALU alu(
		.io_fn(alu_io_fn),
		.io_in2(alu_io_in2),
		.io_in1(alu_io_in1),
		.io_out(alu_io_out),
		.io_adder_out(alu_io_adder_out),
		.io_cmp_out(alu_io_cmp_out)
	);
	MulDiv div(
		.clock(div_clock),
		.reset(div_reset),
		.io_req_ready(div_io_req_ready),
		.io_req_valid(div_io_req_valid),
		.io_req_bits_fn(div_io_req_bits_fn),
		.io_req_bits_in1(div_io_req_bits_in1),
		.io_req_bits_in2(div_io_req_bits_in2),
		.io_req_bits_tag(div_io_req_bits_tag),
		.io_kill(div_io_kill),
		.io_resp_ready(div_io_resp_ready),
		.io_resp_valid(div_io_resp_valid),
		.io_resp_bits_data(div_io_resp_bits_data),
		.io_resp_bits_tag(div_io_resp_bits_tag)
	);
	PlusArgTimeout PlusArgTimeout(
		.clock(PlusArgTimeout_clock),
		.reset(PlusArgTimeout_reset),
		.io_count(PlusArgTimeout_io_count)
	);
	assign rf_id_rs_MPORT_en = 1'h1;
	assign rf_id_rs_MPORT_addr = ~id_raddr1;
	assign rf_id_rs_MPORT_data = rf[rf_id_rs_MPORT_addr];
	assign rf_id_rs_MPORT_1_en = 1'h1;
	assign rf_id_rs_MPORT_1_addr = ~id_raddr2;
	assign rf_id_rs_MPORT_1_data = rf[rf_id_rs_MPORT_1_addr];
	assign rf_MPORT_data = (_rf_wdata_T ? io_dmem_resp_bits_data : _rf_wdata_T_5);
	assign rf_MPORT_addr = ~rf_waddr;
	assign rf_MPORT_mask = 1'h1;
	assign rf_MPORT_en = rf_wen & _T_129;
	assign io_imem_might_request = imem_might_request_reg;
	assign io_imem_req_valid = take_pc_wb | take_pc_mem;
	assign io_imem_req_bits_pc = (wb_xcpt | csr_io_eret ? csr_io_evec : _io_imem_req_bits_pc_T_1);
	assign io_imem_req_bits_speculative = ~take_pc_wb;
	assign io_imem_resp_ready = ibuf_io_imem_ready;
	assign io_imem_btb_update_valid = ((mem_reg_valid & _wb_reg_replay_T) & mem_wrong_npc) & (~mem_cfi | mem_cfi_taken);
	assign io_imem_bht_update_valid = mem_reg_valid & _wb_reg_replay_T;
	assign io_imem_flush_icache = (wb_reg_valid & wb_ctrl_fence_i) & ~io_dmem_s2_nack;
	assign io_dmem_req_valid = ex_reg_valid & ex_ctrl_mem;
	assign io_dmem_req_bits_addr = alu_io_adder_out;
	assign io_dmem_req_bits_tag = {1'd0, ex_dcache_tag};
	assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
	assign io_dmem_req_bits_size = ex_reg_mem_size;
	assign io_dmem_req_bits_signed = ~ex_reg_inst[14];
	assign io_dmem_req_bits_dv = 1'h0;
	assign io_dmem_s1_kill = killm_common | mem_ldst_xcpt;
	assign io_dmem_s1_data_data = mem_reg_rs2;
	assign io_ptw_status_debug = csr_io_status_debug;
	assign io_ptw_pmp_0_cfg_l = csr_io_pmp_0_cfg_l;
	assign io_ptw_pmp_0_cfg_a = csr_io_pmp_0_cfg_a;
	assign io_ptw_pmp_0_cfg_x = csr_io_pmp_0_cfg_x;
	assign io_ptw_pmp_0_cfg_w = csr_io_pmp_0_cfg_w;
	assign io_ptw_pmp_0_cfg_r = csr_io_pmp_0_cfg_r;
	assign io_ptw_pmp_0_addr = csr_io_pmp_0_addr;
	assign io_ptw_pmp_0_mask = csr_io_pmp_0_mask;
	assign io_ptw_pmp_1_cfg_l = csr_io_pmp_1_cfg_l;
	assign io_ptw_pmp_1_cfg_a = csr_io_pmp_1_cfg_a;
	assign io_ptw_pmp_1_cfg_x = csr_io_pmp_1_cfg_x;
	assign io_ptw_pmp_1_cfg_w = csr_io_pmp_1_cfg_w;
	assign io_ptw_pmp_1_cfg_r = csr_io_pmp_1_cfg_r;
	assign io_ptw_pmp_1_addr = csr_io_pmp_1_addr;
	assign io_ptw_pmp_1_mask = csr_io_pmp_1_mask;
	assign io_ptw_pmp_2_cfg_l = csr_io_pmp_2_cfg_l;
	assign io_ptw_pmp_2_cfg_a = csr_io_pmp_2_cfg_a;
	assign io_ptw_pmp_2_cfg_x = csr_io_pmp_2_cfg_x;
	assign io_ptw_pmp_2_cfg_w = csr_io_pmp_2_cfg_w;
	assign io_ptw_pmp_2_cfg_r = csr_io_pmp_2_cfg_r;
	assign io_ptw_pmp_2_addr = csr_io_pmp_2_addr;
	assign io_ptw_pmp_2_mask = csr_io_pmp_2_mask;
	assign io_ptw_pmp_3_cfg_l = csr_io_pmp_3_cfg_l;
	assign io_ptw_pmp_3_cfg_a = csr_io_pmp_3_cfg_a;
	assign io_ptw_pmp_3_cfg_x = csr_io_pmp_3_cfg_x;
	assign io_ptw_pmp_3_cfg_w = csr_io_pmp_3_cfg_w;
	assign io_ptw_pmp_3_cfg_r = csr_io_pmp_3_cfg_r;
	assign io_ptw_pmp_3_addr = csr_io_pmp_3_addr;
	assign io_ptw_pmp_3_mask = csr_io_pmp_3_mask;
	assign io_ptw_pmp_4_cfg_l = csr_io_pmp_4_cfg_l;
	assign io_ptw_pmp_4_cfg_a = csr_io_pmp_4_cfg_a;
	assign io_ptw_pmp_4_cfg_x = csr_io_pmp_4_cfg_x;
	assign io_ptw_pmp_4_cfg_w = csr_io_pmp_4_cfg_w;
	assign io_ptw_pmp_4_cfg_r = csr_io_pmp_4_cfg_r;
	assign io_ptw_pmp_4_addr = csr_io_pmp_4_addr;
	assign io_ptw_pmp_4_mask = csr_io_pmp_4_mask;
	assign io_ptw_pmp_5_cfg_l = csr_io_pmp_5_cfg_l;
	assign io_ptw_pmp_5_cfg_a = csr_io_pmp_5_cfg_a;
	assign io_ptw_pmp_5_cfg_x = csr_io_pmp_5_cfg_x;
	assign io_ptw_pmp_5_cfg_w = csr_io_pmp_5_cfg_w;
	assign io_ptw_pmp_5_cfg_r = csr_io_pmp_5_cfg_r;
	assign io_ptw_pmp_5_addr = csr_io_pmp_5_addr;
	assign io_ptw_pmp_5_mask = csr_io_pmp_5_mask;
	assign io_ptw_pmp_6_cfg_l = csr_io_pmp_6_cfg_l;
	assign io_ptw_pmp_6_cfg_a = csr_io_pmp_6_cfg_a;
	assign io_ptw_pmp_6_cfg_x = csr_io_pmp_6_cfg_x;
	assign io_ptw_pmp_6_cfg_w = csr_io_pmp_6_cfg_w;
	assign io_ptw_pmp_6_cfg_r = csr_io_pmp_6_cfg_r;
	assign io_ptw_pmp_6_addr = csr_io_pmp_6_addr;
	assign io_ptw_pmp_6_mask = csr_io_pmp_6_mask;
	assign io_ptw_pmp_7_cfg_l = csr_io_pmp_7_cfg_l;
	assign io_ptw_pmp_7_cfg_a = csr_io_pmp_7_cfg_a;
	assign io_ptw_pmp_7_cfg_x = csr_io_pmp_7_cfg_x;
	assign io_ptw_pmp_7_cfg_w = csr_io_pmp_7_cfg_w;
	assign io_ptw_pmp_7_cfg_r = csr_io_pmp_7_cfg_r;
	assign io_ptw_pmp_7_addr = csr_io_pmp_7_addr;
	assign io_ptw_pmp_7_mask = csr_io_pmp_7_mask;
	assign io_ptw_customCSRs_csrs_0_value = csr_io_customCSRs_0_value;
	assign io_wfi = csr_io_status_wfi;
	assign ibuf_clock = clock;
	assign ibuf_reset = reset;
	assign ibuf_io_imem_valid = io_imem_resp_valid;
	assign ibuf_io_imem_bits_pc = io_imem_resp_bits_pc;
	assign ibuf_io_imem_bits_data = io_imem_resp_bits_data;
	assign ibuf_io_imem_bits_xcpt_ae_inst = io_imem_resp_bits_xcpt_ae_inst;
	assign ibuf_io_imem_bits_replay = io_imem_resp_bits_replay;
	assign ibuf_io_kill = take_pc_wb | take_pc_mem;
	assign ibuf_io_inst_0_ready = ~ctrl_stalld;
	assign csr_clock = clock;
	assign csr_reset = reset;
	assign csr_io_ungated_clock = clock;
	assign csr_io_interrupts_debug = io_interrupts_debug;
	assign csr_io_interrupts_mtip = io_interrupts_mtip;
	assign csr_io_interrupts_msip = io_interrupts_msip;
	assign csr_io_interrupts_meip = io_interrupts_meip;
	assign csr_io_hartid = io_hartid;
	assign csr_io_rw_addr = wb_reg_inst[31:20];
	assign csr_io_rw_cmd = wb_ctrl_csr & _csr_io_rw_cmd_T_1;
	assign csr_io_rw_wdata = wb_reg_wdata;
	assign csr_io_decode_0_inst = ibuf_io_inst_0_bits_inst_bits;
	assign csr_io_exception = (((((wb_reg_xcpt | _T_91) | _T_93) | _T_99) | _T_101) | _T_103) | _T_105;
	assign csr_io_retire = (wb_reg_valid & ~replay_wb_common) & ~wb_xcpt;
	assign csr_io_cause = (wb_reg_xcpt ? wb_reg_cause : {27'd0, _T_119});
	assign csr_io_pc = wb_reg_pc;
	assign csr_io_tval = (tval_valid ? wb_reg_wdata : 32'h00000000);
	assign csr_io_gva = wb_xcpt & (tval_dmem_addr & wb_reg_hls_or_dv);
	assign csr_io_inst_0 = {_csr_io_inst_0_T_3, wb_reg_raw_inst[15:0]};
	assign bpu_io_status_debug = csr_io_status_debug;
	assign bpu_io_bp_0_control_action = csr_io_bp_0_control_action;
	assign bpu_io_bp_0_control_tmatch = csr_io_bp_0_control_tmatch;
	assign bpu_io_bp_0_control_x = csr_io_bp_0_control_x;
	assign bpu_io_bp_0_control_w = csr_io_bp_0_control_w;
	assign bpu_io_bp_0_control_r = csr_io_bp_0_control_r;
	assign bpu_io_bp_0_address = csr_io_bp_0_address;
	assign bpu_io_pc = ibuf_io_pc;
	assign bpu_io_ea = mem_reg_wdata;
	assign alu_io_fn = ex_ctrl_alu_fn;
	assign alu_io_in2 = (2'h1 == ex_ctrl_sel_alu2 ? $signed({{28 {_ex_op2_T_1[3]}}, _ex_op2_T_1}) : $signed(_ex_op2_T_5));
	assign alu_io_in1 = (2'h2 == ex_ctrl_sel_alu1 ? $signed(ex_reg_pc) : $signed(_ex_op1_T_3));
	assign div_clock = clock;
	assign div_reset = reset;
	assign div_io_req_valid = ex_reg_valid & ex_ctrl_div;
	assign div_io_req_bits_fn = ex_ctrl_alu_fn;
	assign div_io_req_bits_in1 = (ex_reg_rs_bypass_0 ? _ex_rs_T_5 : _ex_rs_T_6);
	assign div_io_req_bits_in2 = (ex_reg_rs_bypass_1 ? _ex_rs_T_12 : _ex_rs_T_13);
	assign div_io_req_bits_tag = ex_reg_inst[11:7];
	assign div_io_kill = killm_common & div_io_kill_REG;
	assign div_io_resp_ready = (dmem_resp_replay & dmem_resp_xpu ? 1'h0 : _ctrl_stalld_T_17);
	assign PlusArgTimeout_clock = clock;
	assign PlusArgTimeout_reset = reset;
	assign PlusArgTimeout_io_count = csr_io_time;
	always @(posedge clock) begin
		if (rf_MPORT_en & rf_MPORT_mask)
			rf[rf_MPORT_addr] <= rf_MPORT_data;
		if (unpause)
			id_reg_pause <= 1'h0;
		else if (_ex_reg_valid_T)
			id_reg_pause <= _GEN_1;
		imem_might_request_reg <= (ex_pc_valid | mem_pc_valid) | io_ptw_customCSRs_csrs_0_value[1];
		if (_ex_reg_valid_T)
			ex_ctrl_branch <= id_ctrl_decoder_3;
		if (_ex_reg_valid_T)
			ex_ctrl_jal <= id_ctrl_decoder_4;
		if (_ex_reg_valid_T)
			ex_ctrl_jalr <= id_ctrl_decoder_5;
		if (_ex_reg_valid_T)
			ex_ctrl_rxs2 <= id_ctrl_decoder_6;
		if (_ex_reg_valid_T)
			ex_ctrl_rxs1 <= id_ctrl_decoder_7;
		if (_ex_reg_valid_T)
			if (id_xcpt) begin
				if (bpu_io_xcpt_if | |_T_37)
					ex_ctrl_sel_alu2 <= 2'h0;
				else if (|_T_35)
					ex_ctrl_sel_alu2 <= 2'h1;
				else
					ex_ctrl_sel_alu2 <= 2'h0;
			end
			else
				ex_ctrl_sel_alu2 <= id_ctrl_decoder_9;
		if (_ex_reg_valid_T)
			if (id_xcpt) begin
				if (bpu_io_xcpt_if | |_T_37)
					ex_ctrl_sel_alu1 <= 2'h2;
				else if (|_T_35)
					ex_ctrl_sel_alu1 <= 2'h2;
				else
					ex_ctrl_sel_alu1 <= 2'h1;
			end
			else
				ex_ctrl_sel_alu1 <= id_ctrl_decoder_10;
		if (_ex_reg_valid_T)
			ex_ctrl_sel_imm <= id_ctrl_decoder_11;
		if (_ex_reg_valid_T)
			if (id_xcpt)
				ex_ctrl_alu_fn <= 4'h0;
			else
				ex_ctrl_alu_fn <= id_ctrl_decoder_13;
		if (_ex_reg_valid_T)
			ex_ctrl_mem <= id_ctrl_decoder_14;
		if (_ex_reg_valid_T)
			ex_ctrl_mem_cmd <= id_ctrl_decoder_15;
		if (_ex_reg_valid_T)
			ex_ctrl_div <= id_ctrl_decoder_21;
		if (_ex_reg_valid_T)
			ex_ctrl_wxd <= id_ctrl_decoder_22;
		if (_ex_reg_valid_T)
			if (id_system_insn & id_ctrl_decoder_14)
				ex_ctrl_csr <= 3'h0;
			else if (id_csr_ren)
				ex_ctrl_csr <= 3'h2;
			else
				ex_ctrl_csr <= id_ctrl_decoder_23;
		if (_ex_reg_valid_T)
			ex_ctrl_fence_i <= id_ctrl_decoder_24;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_ctrl_branch <= ex_ctrl_branch;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_ctrl_jal <= ex_ctrl_jal;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_ctrl_jalr <= ex_ctrl_jalr;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_ctrl_rxs2 <= ex_ctrl_rxs2;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_ctrl_rxs1 <= ex_ctrl_rxs1;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_ctrl_mem <= ex_ctrl_mem;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_ctrl_div <= ex_ctrl_div;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_ctrl_wxd <= ex_ctrl_wxd;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_ctrl_csr <= ex_ctrl_csr;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_ctrl_fence_i <= _GEN_79;
		if (mem_pc_valid)
			wb_ctrl_rxs2 <= mem_ctrl_rxs2;
		if (mem_pc_valid)
			wb_ctrl_rxs1 <= mem_ctrl_rxs1;
		if (mem_pc_valid)
			wb_ctrl_mem <= mem_ctrl_mem;
		if (mem_pc_valid)
			wb_ctrl_div <= mem_ctrl_div;
		if (mem_pc_valid)
			wb_ctrl_wxd <= mem_ctrl_wxd;
		if (mem_pc_valid)
			wb_ctrl_csr <= mem_ctrl_csr;
		if (mem_pc_valid)
			wb_ctrl_fence_i <= mem_ctrl_fence_i;
		ex_reg_xcpt_interrupt <= _ex_reg_replay_T_1 & csr_io_interrupt;
		ex_reg_valid <= ~ctrl_killd;
		if (_ex_reg_valid_T)
			if (id_xcpt)
				ex_reg_rvc <= _GEN_5;
			else
				ex_reg_rvc <= ibuf_io_inst_0_bits_rvc;
		ex_reg_xcpt <= _ex_reg_valid_T & id_xcpt;
		if (_ex_reg_valid_T)
			ex_reg_flush_pipe <= id_ctrl_decoder_24 | id_csr_flush;
		if (_ex_reg_valid_T)
			ex_reg_load_use <= id_load_use;
		if ((_ex_reg_valid_T | csr_io_interrupt) | ibuf_io_inst_0_bits_replay)
			if (csr_io_interrupt)
				ex_reg_cause <= csr_io_interrupt_cause;
			else
				ex_reg_cause <= {27'd0, _T_18};
		ex_reg_replay <= (~take_pc_mem_wb & ibuf_io_inst_0_valid) & ibuf_io_inst_0_bits_replay;
		if ((_ex_reg_valid_T | csr_io_interrupt) | ibuf_io_inst_0_bits_replay)
			ex_reg_pc <= ibuf_io_pc;
		if (_ex_reg_valid_T)
			if (_T_46)
				ex_reg_mem_size <= _ex_reg_mem_size_T_6;
			else
				ex_reg_mem_size <= ibuf_io_inst_0_bits_inst_bits[13:12];
		if ((_ex_reg_valid_T | csr_io_interrupt) | ibuf_io_inst_0_bits_replay)
			ex_reg_inst <= ibuf_io_inst_0_bits_inst_bits;
		if ((_ex_reg_valid_T | csr_io_interrupt) | ibuf_io_inst_0_bits_replay)
			ex_reg_raw_inst <= ibuf_io_inst_0_bits_raw;
		mem_reg_xcpt_interrupt <= _ex_reg_replay_T & ex_reg_xcpt_interrupt;
		mem_reg_valid <= ~ctrl_killx;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_reg_rvc <= ex_reg_rvc;
		mem_reg_xcpt <= _mem_reg_valid_T & ex_xcpt;
		mem_reg_replay <= _ex_reg_replay_T & replay_ex;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_reg_flush_pipe <= _GEN_80;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_reg_cause <= ex_reg_cause;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_reg_slow_bypass <= ex_slow_bypass;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_reg_load <= ex_ctrl_mem & _mem_reg_load_T_24;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_reg_store <= ex_ctrl_mem & _mem_reg_store_T_22;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_reg_pc <= ex_reg_pc;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_reg_inst <= ex_reg_inst;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_reg_hls_or_dv <= io_dmem_req_bits_dv;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_reg_raw_inst <= ex_reg_raw_inst;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_reg_wdata <= _mem_reg_wdata_T;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				if (ex_ctrl_rxs2 & ex_ctrl_mem)
					if (ex_reg_mem_size == 2'h0)
						mem_reg_rs2 <= _mem_reg_rs2_T_3;
					else
						mem_reg_rs2 <= _mem_reg_rs2_T_7;
		if (!(mem_reg_valid & mem_reg_flush_pipe))
			if (ex_pc_valid)
				mem_br_taken <= alu_io_cmp_out;
		wb_reg_valid <= ~ctrl_killm;
		wb_reg_xcpt <= mem_xcpt & _wb_reg_replay_T;
		wb_reg_replay <= replay_mem & ~take_pc_wb;
		wb_reg_flush_pipe <= _wb_reg_valid_T & mem_reg_flush_pipe;
		if (mem_pc_valid)
			if (_T_70)
				wb_reg_cause <= mem_reg_cause;
			else
				wb_reg_cause <= {28'd0, _T_74};
		if (mem_pc_valid)
			wb_reg_pc <= mem_reg_pc;
		if (mem_pc_valid)
			wb_reg_hls_or_dv <= mem_reg_hls_or_dv;
		if (mem_pc_valid)
			wb_reg_inst <= mem_reg_inst;
		if (mem_pc_valid)
			wb_reg_raw_inst <= mem_reg_raw_inst;
		if (mem_pc_valid)
			wb_reg_wdata <= mem_int_wdata;
		if (reset)
			id_reg_fence <= 1'h0;
		else if (_ex_reg_valid_T)
			id_reg_fence <= _GEN_2;
		else if (~id_mem_busy)
			id_reg_fence <= 1'h0;
		if (_ex_reg_valid_T)
			if (id_illegal_insn)
				ex_reg_rs_bypass_0 <= 1'h0;
			else
				ex_reg_rs_bypass_0 <= do_bypass;
		if (_ex_reg_valid_T)
			ex_reg_rs_bypass_1 <= do_bypass_1;
		if (_ex_reg_valid_T)
			if (id_illegal_insn)
				ex_reg_rs_lsb_0 <= inst[1:0];
			else if (id_ctrl_decoder_7 & ~do_bypass)
				ex_reg_rs_lsb_0 <= id_rs_0[1:0];
			else if (id_bypass_src_0_0)
				ex_reg_rs_lsb_0 <= 2'h0;
			else
				ex_reg_rs_lsb_0 <= _bypass_src_T_1;
		if (_ex_reg_valid_T)
			if (id_ctrl_decoder_6 & ~do_bypass_1)
				ex_reg_rs_lsb_1 <= id_rs_1[1:0];
			else if (id_bypass_src_1_0)
				ex_reg_rs_lsb_1 <= 2'h0;
			else if (id_bypass_src_1_1)
				ex_reg_rs_lsb_1 <= 2'h1;
			else
				ex_reg_rs_lsb_1 <= _bypass_src_T_2;
		if (_ex_reg_valid_T)
			if (id_illegal_insn)
				ex_reg_rs_msb_0 <= inst[31:2];
			else if (id_ctrl_decoder_7 & ~do_bypass)
				ex_reg_rs_msb_0 <= id_rs_0[31:2];
		if (_ex_reg_valid_T)
			if (id_ctrl_decoder_6 & ~do_bypass_1)
				ex_reg_rs_msb_1 <= id_rs_1[31:2];
		if (reset)
			_r <= 32'h00000000;
		else if (_T_149)
			_r <= _T_148;
		else if (ll_wen)
			_r <= _T_143;
		blocked <= (_replay_ex_structural_T & _dcache_blocked_T) & ((blocked | io_dmem_req_valid) | io_dmem_s2_nack);
		div_io_kill_REG <= div_io_req_ready & div_io_req_valid;
		if (ex_reg_rs_bypass_0) begin
			if (ex_reg_rs_lsb_0 == 2'h3)
				coreMonitorBundle_rd0val_x23 <= io_dmem_resp_bits_data_word_bypass;
			else if (ex_reg_rs_lsb_0 == 2'h2)
				coreMonitorBundle_rd0val_x23 <= wb_reg_wdata;
			else if (ex_reg_rs_lsb_0 == 2'h1)
				coreMonitorBundle_rd0val_x23 <= mem_reg_wdata;
			else
				coreMonitorBundle_rd0val_x23 <= 32'h00000000;
		end
		else
			coreMonitorBundle_rd0val_x23 <= _ex_rs_T_6;
		coreMonitorBundle_rd0val_REG <= coreMonitorBundle_rd0val_x23;
		if (ex_reg_rs_bypass_1) begin
			if (ex_reg_rs_lsb_1 == 2'h3)
				coreMonitorBundle_rd1val_x29 <= io_dmem_resp_bits_data_word_bypass;
			else if (ex_reg_rs_lsb_1 == 2'h2)
				coreMonitorBundle_rd1val_x29 <= wb_reg_wdata;
			else if (ex_reg_rs_lsb_1 == 2'h1)
				coreMonitorBundle_rd1val_x29 <= mem_reg_wdata;
			else
				coreMonitorBundle_rd1val_x29 <= 32'h00000000;
		end
		else
			coreMonitorBundle_rd1val_x29 <= _ex_rs_T_13;
		coreMonitorBundle_rd1val_REG <= coreMonitorBundle_rd1val_x29;
	end
endmodule
module RocketTile (
	clock,
	reset,
	auto_slave_in_a_ready,
	auto_slave_in_a_valid,
	auto_slave_in_a_bits_opcode,
	auto_slave_in_a_bits_param,
	auto_slave_in_a_bits_size,
	auto_slave_in_a_bits_source,
	auto_slave_in_a_bits_address,
	auto_slave_in_a_bits_mask,
	auto_slave_in_a_bits_data,
	auto_slave_in_d_ready,
	auto_slave_in_d_valid,
	auto_slave_in_d_bits_opcode,
	auto_slave_in_d_bits_size,
	auto_slave_in_d_bits_source,
	auto_slave_in_d_bits_data,
	auto_wfi_out_0,
	auto_int_local_in_2_0,
	auto_int_local_in_1_0,
	auto_int_local_in_1_1,
	auto_int_local_in_0_0,
	auto_hartid_in,
	auto_tl_other_masters_out_a_ready,
	auto_tl_other_masters_out_a_valid,
	auto_tl_other_masters_out_a_bits_opcode,
	auto_tl_other_masters_out_a_bits_param,
	auto_tl_other_masters_out_a_bits_size,
	auto_tl_other_masters_out_a_bits_source,
	auto_tl_other_masters_out_a_bits_address,
	auto_tl_other_masters_out_a_bits_mask,
	auto_tl_other_masters_out_a_bits_data,
	auto_tl_other_masters_out_d_ready,
	auto_tl_other_masters_out_d_valid,
	auto_tl_other_masters_out_d_bits_opcode,
	auto_tl_other_masters_out_d_bits_param,
	auto_tl_other_masters_out_d_bits_size,
	auto_tl_other_masters_out_d_bits_source,
	auto_tl_other_masters_out_d_bits_sink,
	auto_tl_other_masters_out_d_bits_denied,
	auto_tl_other_masters_out_d_bits_data,
	auto_tl_other_masters_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_slave_in_a_ready;
	input auto_slave_in_a_valid;
	input [2:0] auto_slave_in_a_bits_opcode;
	input [2:0] auto_slave_in_a_bits_param;
	input [2:0] auto_slave_in_a_bits_size;
	input [2:0] auto_slave_in_a_bits_source;
	input [31:0] auto_slave_in_a_bits_address;
	input [3:0] auto_slave_in_a_bits_mask;
	input [31:0] auto_slave_in_a_bits_data;
	input auto_slave_in_d_ready;
	output wire auto_slave_in_d_valid;
	output wire [2:0] auto_slave_in_d_bits_opcode;
	output wire [2:0] auto_slave_in_d_bits_size;
	output wire [2:0] auto_slave_in_d_bits_source;
	output wire [31:0] auto_slave_in_d_bits_data;
	output wire auto_wfi_out_0;
	input auto_int_local_in_2_0;
	input auto_int_local_in_1_0;
	input auto_int_local_in_1_1;
	input auto_int_local_in_0_0;
	input auto_hartid_in;
	input auto_tl_other_masters_out_a_ready;
	output wire auto_tl_other_masters_out_a_valid;
	output wire [2:0] auto_tl_other_masters_out_a_bits_opcode;
	output wire [2:0] auto_tl_other_masters_out_a_bits_param;
	output wire [3:0] auto_tl_other_masters_out_a_bits_size;
	output wire auto_tl_other_masters_out_a_bits_source;
	output wire [31:0] auto_tl_other_masters_out_a_bits_address;
	output wire [3:0] auto_tl_other_masters_out_a_bits_mask;
	output wire [31:0] auto_tl_other_masters_out_a_bits_data;
	output wire auto_tl_other_masters_out_d_ready;
	input auto_tl_other_masters_out_d_valid;
	input [2:0] auto_tl_other_masters_out_d_bits_opcode;
	input [1:0] auto_tl_other_masters_out_d_bits_param;
	input [3:0] auto_tl_other_masters_out_d_bits_size;
	input auto_tl_other_masters_out_d_bits_source;
	input auto_tl_other_masters_out_d_bits_sink;
	input auto_tl_other_masters_out_d_bits_denied;
	input [31:0] auto_tl_other_masters_out_d_bits_data;
	input auto_tl_other_masters_out_d_bits_corrupt;
	wire tlMasterXbar_clock;
	wire tlMasterXbar_reset;
	wire tlMasterXbar_auto_in_1_a_ready;
	wire tlMasterXbar_auto_in_1_a_valid;
	wire [31:0] tlMasterXbar_auto_in_1_a_bits_address;
	wire tlMasterXbar_auto_in_1_d_valid;
	wire [2:0] tlMasterXbar_auto_in_1_d_bits_opcode;
	wire [3:0] tlMasterXbar_auto_in_1_d_bits_size;
	wire [31:0] tlMasterXbar_auto_in_1_d_bits_data;
	wire tlMasterXbar_auto_in_1_d_bits_corrupt;
	wire tlMasterXbar_auto_in_0_a_ready;
	wire tlMasterXbar_auto_in_0_a_valid;
	wire [2:0] tlMasterXbar_auto_in_0_a_bits_opcode;
	wire [2:0] tlMasterXbar_auto_in_0_a_bits_param;
	wire [3:0] tlMasterXbar_auto_in_0_a_bits_size;
	wire [31:0] tlMasterXbar_auto_in_0_a_bits_address;
	wire [3:0] tlMasterXbar_auto_in_0_a_bits_mask;
	wire [31:0] tlMasterXbar_auto_in_0_a_bits_data;
	wire tlMasterXbar_auto_in_0_d_ready;
	wire tlMasterXbar_auto_in_0_d_valid;
	wire [2:0] tlMasterXbar_auto_in_0_d_bits_opcode;
	wire [3:0] tlMasterXbar_auto_in_0_d_bits_size;
	wire tlMasterXbar_auto_in_0_d_bits_denied;
	wire [31:0] tlMasterXbar_auto_in_0_d_bits_data;
	wire tlMasterXbar_auto_out_a_ready;
	wire tlMasterXbar_auto_out_a_valid;
	wire [2:0] tlMasterXbar_auto_out_a_bits_opcode;
	wire [2:0] tlMasterXbar_auto_out_a_bits_param;
	wire [3:0] tlMasterXbar_auto_out_a_bits_size;
	wire tlMasterXbar_auto_out_a_bits_source;
	wire [31:0] tlMasterXbar_auto_out_a_bits_address;
	wire [3:0] tlMasterXbar_auto_out_a_bits_mask;
	wire [31:0] tlMasterXbar_auto_out_a_bits_data;
	wire tlMasterXbar_auto_out_d_ready;
	wire tlMasterXbar_auto_out_d_valid;
	wire [2:0] tlMasterXbar_auto_out_d_bits_opcode;
	wire [1:0] tlMasterXbar_auto_out_d_bits_param;
	wire [3:0] tlMasterXbar_auto_out_d_bits_size;
	wire tlMasterXbar_auto_out_d_bits_source;
	wire tlMasterXbar_auto_out_d_bits_sink;
	wire tlMasterXbar_auto_out_d_bits_denied;
	wire [31:0] tlMasterXbar_auto_out_d_bits_data;
	wire tlMasterXbar_auto_out_d_bits_corrupt;
	wire tlSlaveXbar_auto_in_a_ready;
	wire tlSlaveXbar_auto_in_a_valid;
	wire [2:0] tlSlaveXbar_auto_in_a_bits_opcode;
	wire [2:0] tlSlaveXbar_auto_in_a_bits_param;
	wire [2:0] tlSlaveXbar_auto_in_a_bits_size;
	wire [2:0] tlSlaveXbar_auto_in_a_bits_source;
	wire [31:0] tlSlaveXbar_auto_in_a_bits_address;
	wire [3:0] tlSlaveXbar_auto_in_a_bits_mask;
	wire [31:0] tlSlaveXbar_auto_in_a_bits_data;
	wire tlSlaveXbar_auto_in_d_ready;
	wire tlSlaveXbar_auto_in_d_valid;
	wire [2:0] tlSlaveXbar_auto_in_d_bits_opcode;
	wire [2:0] tlSlaveXbar_auto_in_d_bits_size;
	wire [2:0] tlSlaveXbar_auto_in_d_bits_source;
	wire [31:0] tlSlaveXbar_auto_in_d_bits_data;
	wire tlSlaveXbar_auto_out_a_ready;
	wire tlSlaveXbar_auto_out_a_valid;
	wire [2:0] tlSlaveXbar_auto_out_a_bits_opcode;
	wire [2:0] tlSlaveXbar_auto_out_a_bits_param;
	wire [2:0] tlSlaveXbar_auto_out_a_bits_size;
	wire [2:0] tlSlaveXbar_auto_out_a_bits_source;
	wire [31:0] tlSlaveXbar_auto_out_a_bits_address;
	wire [3:0] tlSlaveXbar_auto_out_a_bits_mask;
	wire [31:0] tlSlaveXbar_auto_out_a_bits_data;
	wire tlSlaveXbar_auto_out_d_ready;
	wire tlSlaveXbar_auto_out_d_valid;
	wire [2:0] tlSlaveXbar_auto_out_d_bits_opcode;
	wire [2:0] tlSlaveXbar_auto_out_d_bits_size;
	wire [2:0] tlSlaveXbar_auto_out_d_bits_source;
	wire [31:0] tlSlaveXbar_auto_out_d_bits_data;
	wire intXbar_auto_int_in_2_0;
	wire intXbar_auto_int_in_1_0;
	wire intXbar_auto_int_in_1_1;
	wire intXbar_auto_int_in_0_0;
	wire intXbar_auto_int_out_0;
	wire intXbar_auto_int_out_1;
	wire intXbar_auto_int_out_2;
	wire intXbar_auto_int_out_3;
	wire broadcast_auto_in;
	wire broadcast_auto_out_0;
	wire dcache_clock;
	wire dcache_reset;
	wire dcache_auto_out_a_ready;
	wire dcache_auto_out_a_valid;
	wire [2:0] dcache_auto_out_a_bits_opcode;
	wire [2:0] dcache_auto_out_a_bits_param;
	wire [3:0] dcache_auto_out_a_bits_size;
	wire [31:0] dcache_auto_out_a_bits_address;
	wire [3:0] dcache_auto_out_a_bits_mask;
	wire [31:0] dcache_auto_out_a_bits_data;
	wire dcache_auto_out_d_ready;
	wire dcache_auto_out_d_valid;
	wire [2:0] dcache_auto_out_d_bits_opcode;
	wire [3:0] dcache_auto_out_d_bits_size;
	wire dcache_auto_out_d_bits_denied;
	wire [31:0] dcache_auto_out_d_bits_data;
	wire dcache_io_cpu_req_ready;
	wire dcache_io_cpu_req_valid;
	wire [31:0] dcache_io_cpu_req_bits_addr;
	wire [6:0] dcache_io_cpu_req_bits_tag;
	wire [4:0] dcache_io_cpu_req_bits_cmd;
	wire [1:0] dcache_io_cpu_req_bits_size;
	wire dcache_io_cpu_req_bits_signed;
	wire [1:0] dcache_io_cpu_req_bits_dprv;
	wire dcache_io_cpu_req_bits_no_xcpt;
	wire dcache_io_cpu_s1_kill;
	wire [31:0] dcache_io_cpu_s1_data_data;
	wire [3:0] dcache_io_cpu_s1_data_mask;
	wire dcache_io_cpu_s2_nack;
	wire dcache_io_cpu_resp_valid;
	wire [31:0] dcache_io_cpu_resp_bits_addr;
	wire [6:0] dcache_io_cpu_resp_bits_tag;
	wire [4:0] dcache_io_cpu_resp_bits_cmd;
	wire [1:0] dcache_io_cpu_resp_bits_size;
	wire dcache_io_cpu_resp_bits_signed;
	wire [1:0] dcache_io_cpu_resp_bits_dprv;
	wire dcache_io_cpu_resp_bits_dv;
	wire [31:0] dcache_io_cpu_resp_bits_data;
	wire [3:0] dcache_io_cpu_resp_bits_mask;
	wire dcache_io_cpu_resp_bits_replay;
	wire dcache_io_cpu_resp_bits_has_data;
	wire [31:0] dcache_io_cpu_resp_bits_data_word_bypass;
	wire [31:0] dcache_io_cpu_resp_bits_data_raw;
	wire [31:0] dcache_io_cpu_resp_bits_store_data;
	wire dcache_io_cpu_replay_next;
	wire dcache_io_cpu_s2_xcpt_ma_ld;
	wire dcache_io_cpu_s2_xcpt_ma_st;
	wire dcache_io_cpu_s2_xcpt_pf_ld;
	wire dcache_io_cpu_s2_xcpt_pf_st;
	wire dcache_io_cpu_s2_xcpt_gf_ld;
	wire dcache_io_cpu_s2_xcpt_gf_st;
	wire dcache_io_cpu_s2_xcpt_ae_ld;
	wire dcache_io_cpu_s2_xcpt_ae_st;
	wire dcache_io_cpu_ordered;
	wire dcache_io_cpu_perf_grant;
	wire dcache_io_ptw_status_debug;
	wire dcache_io_ptw_pmp_0_cfg_l;
	wire [1:0] dcache_io_ptw_pmp_0_cfg_a;
	wire dcache_io_ptw_pmp_0_cfg_x;
	wire dcache_io_ptw_pmp_0_cfg_w;
	wire dcache_io_ptw_pmp_0_cfg_r;
	wire [29:0] dcache_io_ptw_pmp_0_addr;
	wire [31:0] dcache_io_ptw_pmp_0_mask;
	wire dcache_io_ptw_pmp_1_cfg_l;
	wire [1:0] dcache_io_ptw_pmp_1_cfg_a;
	wire dcache_io_ptw_pmp_1_cfg_x;
	wire dcache_io_ptw_pmp_1_cfg_w;
	wire dcache_io_ptw_pmp_1_cfg_r;
	wire [29:0] dcache_io_ptw_pmp_1_addr;
	wire [31:0] dcache_io_ptw_pmp_1_mask;
	wire dcache_io_ptw_pmp_2_cfg_l;
	wire [1:0] dcache_io_ptw_pmp_2_cfg_a;
	wire dcache_io_ptw_pmp_2_cfg_x;
	wire dcache_io_ptw_pmp_2_cfg_w;
	wire dcache_io_ptw_pmp_2_cfg_r;
	wire [29:0] dcache_io_ptw_pmp_2_addr;
	wire [31:0] dcache_io_ptw_pmp_2_mask;
	wire dcache_io_ptw_pmp_3_cfg_l;
	wire [1:0] dcache_io_ptw_pmp_3_cfg_a;
	wire dcache_io_ptw_pmp_3_cfg_x;
	wire dcache_io_ptw_pmp_3_cfg_w;
	wire dcache_io_ptw_pmp_3_cfg_r;
	wire [29:0] dcache_io_ptw_pmp_3_addr;
	wire [31:0] dcache_io_ptw_pmp_3_mask;
	wire dcache_io_ptw_pmp_4_cfg_l;
	wire [1:0] dcache_io_ptw_pmp_4_cfg_a;
	wire dcache_io_ptw_pmp_4_cfg_x;
	wire dcache_io_ptw_pmp_4_cfg_w;
	wire dcache_io_ptw_pmp_4_cfg_r;
	wire [29:0] dcache_io_ptw_pmp_4_addr;
	wire [31:0] dcache_io_ptw_pmp_4_mask;
	wire dcache_io_ptw_pmp_5_cfg_l;
	wire [1:0] dcache_io_ptw_pmp_5_cfg_a;
	wire dcache_io_ptw_pmp_5_cfg_x;
	wire dcache_io_ptw_pmp_5_cfg_w;
	wire dcache_io_ptw_pmp_5_cfg_r;
	wire [29:0] dcache_io_ptw_pmp_5_addr;
	wire [31:0] dcache_io_ptw_pmp_5_mask;
	wire dcache_io_ptw_pmp_6_cfg_l;
	wire [1:0] dcache_io_ptw_pmp_6_cfg_a;
	wire dcache_io_ptw_pmp_6_cfg_x;
	wire dcache_io_ptw_pmp_6_cfg_w;
	wire dcache_io_ptw_pmp_6_cfg_r;
	wire [29:0] dcache_io_ptw_pmp_6_addr;
	wire [31:0] dcache_io_ptw_pmp_6_mask;
	wire dcache_io_ptw_pmp_7_cfg_l;
	wire [1:0] dcache_io_ptw_pmp_7_cfg_a;
	wire dcache_io_ptw_pmp_7_cfg_x;
	wire dcache_io_ptw_pmp_7_cfg_w;
	wire dcache_io_ptw_pmp_7_cfg_r;
	wire [29:0] dcache_io_ptw_pmp_7_addr;
	wire [31:0] dcache_io_ptw_pmp_7_mask;
	wire frontend_clock;
	wire frontend_reset;
	wire frontend_auto_icache_master_out_a_ready;
	wire frontend_auto_icache_master_out_a_valid;
	wire [31:0] frontend_auto_icache_master_out_a_bits_address;
	wire frontend_auto_icache_master_out_d_valid;
	wire [2:0] frontend_auto_icache_master_out_d_bits_opcode;
	wire [3:0] frontend_auto_icache_master_out_d_bits_size;
	wire [31:0] frontend_auto_icache_master_out_d_bits_data;
	wire frontend_auto_icache_master_out_d_bits_corrupt;
	wire frontend_io_cpu_might_request;
	wire frontend_io_cpu_req_valid;
	wire [31:0] frontend_io_cpu_req_bits_pc;
	wire frontend_io_cpu_req_bits_speculative;
	wire frontend_io_cpu_resp_ready;
	wire frontend_io_cpu_resp_valid;
	wire [31:0] frontend_io_cpu_resp_bits_pc;
	wire [31:0] frontend_io_cpu_resp_bits_data;
	wire frontend_io_cpu_resp_bits_xcpt_ae_inst;
	wire frontend_io_cpu_resp_bits_replay;
	wire frontend_io_cpu_btb_update_valid;
	wire frontend_io_cpu_bht_update_valid;
	wire frontend_io_cpu_flush_icache;
	wire [31:0] frontend_io_cpu_npc;
	wire frontend_io_ptw_status_debug;
	wire frontend_io_ptw_pmp_0_cfg_l;
	wire [1:0] frontend_io_ptw_pmp_0_cfg_a;
	wire frontend_io_ptw_pmp_0_cfg_x;
	wire frontend_io_ptw_pmp_0_cfg_w;
	wire frontend_io_ptw_pmp_0_cfg_r;
	wire [29:0] frontend_io_ptw_pmp_0_addr;
	wire [31:0] frontend_io_ptw_pmp_0_mask;
	wire frontend_io_ptw_pmp_1_cfg_l;
	wire [1:0] frontend_io_ptw_pmp_1_cfg_a;
	wire frontend_io_ptw_pmp_1_cfg_x;
	wire frontend_io_ptw_pmp_1_cfg_w;
	wire frontend_io_ptw_pmp_1_cfg_r;
	wire [29:0] frontend_io_ptw_pmp_1_addr;
	wire [31:0] frontend_io_ptw_pmp_1_mask;
	wire frontend_io_ptw_pmp_2_cfg_l;
	wire [1:0] frontend_io_ptw_pmp_2_cfg_a;
	wire frontend_io_ptw_pmp_2_cfg_x;
	wire frontend_io_ptw_pmp_2_cfg_w;
	wire frontend_io_ptw_pmp_2_cfg_r;
	wire [29:0] frontend_io_ptw_pmp_2_addr;
	wire [31:0] frontend_io_ptw_pmp_2_mask;
	wire frontend_io_ptw_pmp_3_cfg_l;
	wire [1:0] frontend_io_ptw_pmp_3_cfg_a;
	wire frontend_io_ptw_pmp_3_cfg_x;
	wire frontend_io_ptw_pmp_3_cfg_w;
	wire frontend_io_ptw_pmp_3_cfg_r;
	wire [29:0] frontend_io_ptw_pmp_3_addr;
	wire [31:0] frontend_io_ptw_pmp_3_mask;
	wire frontend_io_ptw_pmp_4_cfg_l;
	wire [1:0] frontend_io_ptw_pmp_4_cfg_a;
	wire frontend_io_ptw_pmp_4_cfg_x;
	wire frontend_io_ptw_pmp_4_cfg_w;
	wire frontend_io_ptw_pmp_4_cfg_r;
	wire [29:0] frontend_io_ptw_pmp_4_addr;
	wire [31:0] frontend_io_ptw_pmp_4_mask;
	wire frontend_io_ptw_pmp_5_cfg_l;
	wire [1:0] frontend_io_ptw_pmp_5_cfg_a;
	wire frontend_io_ptw_pmp_5_cfg_x;
	wire frontend_io_ptw_pmp_5_cfg_w;
	wire frontend_io_ptw_pmp_5_cfg_r;
	wire [29:0] frontend_io_ptw_pmp_5_addr;
	wire [31:0] frontend_io_ptw_pmp_5_mask;
	wire frontend_io_ptw_pmp_6_cfg_l;
	wire [1:0] frontend_io_ptw_pmp_6_cfg_a;
	wire frontend_io_ptw_pmp_6_cfg_x;
	wire frontend_io_ptw_pmp_6_cfg_w;
	wire frontend_io_ptw_pmp_6_cfg_r;
	wire [29:0] frontend_io_ptw_pmp_6_addr;
	wire [31:0] frontend_io_ptw_pmp_6_mask;
	wire frontend_io_ptw_pmp_7_cfg_l;
	wire [1:0] frontend_io_ptw_pmp_7_cfg_a;
	wire frontend_io_ptw_pmp_7_cfg_x;
	wire frontend_io_ptw_pmp_7_cfg_w;
	wire frontend_io_ptw_pmp_7_cfg_r;
	wire [29:0] frontend_io_ptw_pmp_7_addr;
	wire [31:0] frontend_io_ptw_pmp_7_mask;
	wire [31:0] frontend_io_ptw_customCSRs_csrs_0_value;
	wire dtim_adapter_clock;
	wire dtim_adapter_reset;
	wire dtim_adapter_auto_in_a_ready;
	wire dtim_adapter_auto_in_a_valid;
	wire [2:0] dtim_adapter_auto_in_a_bits_opcode;
	wire [2:0] dtim_adapter_auto_in_a_bits_param;
	wire [1:0] dtim_adapter_auto_in_a_bits_size;
	wire [8:0] dtim_adapter_auto_in_a_bits_source;
	wire [31:0] dtim_adapter_auto_in_a_bits_address;
	wire [3:0] dtim_adapter_auto_in_a_bits_mask;
	wire [31:0] dtim_adapter_auto_in_a_bits_data;
	wire dtim_adapter_auto_in_d_ready;
	wire dtim_adapter_auto_in_d_valid;
	wire [2:0] dtim_adapter_auto_in_d_bits_opcode;
	wire [1:0] dtim_adapter_auto_in_d_bits_size;
	wire [8:0] dtim_adapter_auto_in_d_bits_source;
	wire [31:0] dtim_adapter_auto_in_d_bits_data;
	wire dtim_adapter_io_dmem_req_ready;
	wire dtim_adapter_io_dmem_req_valid;
	wire [31:0] dtim_adapter_io_dmem_req_bits_addr;
	wire [4:0] dtim_adapter_io_dmem_req_bits_cmd;
	wire [1:0] dtim_adapter_io_dmem_req_bits_size;
	wire dtim_adapter_io_dmem_s1_kill;
	wire [31:0] dtim_adapter_io_dmem_s1_data_data;
	wire [3:0] dtim_adapter_io_dmem_s1_data_mask;
	wire dtim_adapter_io_dmem_s2_nack;
	wire dtim_adapter_io_dmem_resp_valid;
	wire [31:0] dtim_adapter_io_dmem_resp_bits_data_raw;
	wire fragmenter_1_clock;
	wire fragmenter_1_reset;
	wire fragmenter_1_auto_in_a_ready;
	wire fragmenter_1_auto_in_a_valid;
	wire [2:0] fragmenter_1_auto_in_a_bits_opcode;
	wire [2:0] fragmenter_1_auto_in_a_bits_param;
	wire [2:0] fragmenter_1_auto_in_a_bits_size;
	wire [2:0] fragmenter_1_auto_in_a_bits_source;
	wire [31:0] fragmenter_1_auto_in_a_bits_address;
	wire [3:0] fragmenter_1_auto_in_a_bits_mask;
	wire [31:0] fragmenter_1_auto_in_a_bits_data;
	wire fragmenter_1_auto_in_d_ready;
	wire fragmenter_1_auto_in_d_valid;
	wire [2:0] fragmenter_1_auto_in_d_bits_opcode;
	wire [2:0] fragmenter_1_auto_in_d_bits_size;
	wire [2:0] fragmenter_1_auto_in_d_bits_source;
	wire [31:0] fragmenter_1_auto_in_d_bits_data;
	wire fragmenter_1_auto_out_a_ready;
	wire fragmenter_1_auto_out_a_valid;
	wire [2:0] fragmenter_1_auto_out_a_bits_opcode;
	wire [2:0] fragmenter_1_auto_out_a_bits_param;
	wire [1:0] fragmenter_1_auto_out_a_bits_size;
	wire [8:0] fragmenter_1_auto_out_a_bits_source;
	wire [31:0] fragmenter_1_auto_out_a_bits_address;
	wire [3:0] fragmenter_1_auto_out_a_bits_mask;
	wire [31:0] fragmenter_1_auto_out_a_bits_data;
	wire fragmenter_1_auto_out_d_ready;
	wire fragmenter_1_auto_out_d_valid;
	wire [2:0] fragmenter_1_auto_out_d_bits_opcode;
	wire [1:0] fragmenter_1_auto_out_d_bits_size;
	wire [8:0] fragmenter_1_auto_out_d_bits_source;
	wire [31:0] fragmenter_1_auto_out_d_bits_data;
	wire dcacheArb_clock;
	wire dcacheArb_io_requestor_0_req_ready;
	wire dcacheArb_io_requestor_0_req_valid;
	wire [31:0] dcacheArb_io_requestor_0_req_bits_addr;
	wire [6:0] dcacheArb_io_requestor_0_req_bits_tag;
	wire [4:0] dcacheArb_io_requestor_0_req_bits_cmd;
	wire [1:0] dcacheArb_io_requestor_0_req_bits_size;
	wire dcacheArb_io_requestor_0_req_bits_signed;
	wire dcacheArb_io_requestor_0_s1_kill;
	wire [31:0] dcacheArb_io_requestor_0_s1_data_data;
	wire dcacheArb_io_requestor_0_s2_nack;
	wire dcacheArb_io_requestor_0_resp_valid;
	wire [6:0] dcacheArb_io_requestor_0_resp_bits_tag;
	wire [31:0] dcacheArb_io_requestor_0_resp_bits_data;
	wire dcacheArb_io_requestor_0_resp_bits_replay;
	wire dcacheArb_io_requestor_0_resp_bits_has_data;
	wire [31:0] dcacheArb_io_requestor_0_resp_bits_data_word_bypass;
	wire dcacheArb_io_requestor_0_replay_next;
	wire dcacheArb_io_requestor_0_s2_xcpt_ma_ld;
	wire dcacheArb_io_requestor_0_s2_xcpt_ma_st;
	wire dcacheArb_io_requestor_0_s2_xcpt_pf_ld;
	wire dcacheArb_io_requestor_0_s2_xcpt_pf_st;
	wire dcacheArb_io_requestor_0_s2_xcpt_ae_ld;
	wire dcacheArb_io_requestor_0_s2_xcpt_ae_st;
	wire dcacheArb_io_requestor_0_ordered;
	wire dcacheArb_io_requestor_0_perf_grant;
	wire dcacheArb_io_requestor_1_req_ready;
	wire dcacheArb_io_requestor_1_req_valid;
	wire [31:0] dcacheArb_io_requestor_1_req_bits_addr;
	wire [4:0] dcacheArb_io_requestor_1_req_bits_cmd;
	wire [1:0] dcacheArb_io_requestor_1_req_bits_size;
	wire dcacheArb_io_requestor_1_s1_kill;
	wire [31:0] dcacheArb_io_requestor_1_s1_data_data;
	wire [3:0] dcacheArb_io_requestor_1_s1_data_mask;
	wire dcacheArb_io_requestor_1_s2_nack;
	wire dcacheArb_io_requestor_1_resp_valid;
	wire [31:0] dcacheArb_io_requestor_1_resp_bits_data_raw;
	wire dcacheArb_io_mem_req_ready;
	wire dcacheArb_io_mem_req_valid;
	wire [31:0] dcacheArb_io_mem_req_bits_addr;
	wire [6:0] dcacheArb_io_mem_req_bits_tag;
	wire [4:0] dcacheArb_io_mem_req_bits_cmd;
	wire [1:0] dcacheArb_io_mem_req_bits_size;
	wire dcacheArb_io_mem_req_bits_signed;
	wire [1:0] dcacheArb_io_mem_req_bits_dprv;
	wire dcacheArb_io_mem_req_bits_no_xcpt;
	wire dcacheArb_io_mem_s1_kill;
	wire [31:0] dcacheArb_io_mem_s1_data_data;
	wire [3:0] dcacheArb_io_mem_s1_data_mask;
	wire dcacheArb_io_mem_s2_nack;
	wire dcacheArb_io_mem_resp_valid;
	wire [6:0] dcacheArb_io_mem_resp_bits_tag;
	wire [31:0] dcacheArb_io_mem_resp_bits_data;
	wire dcacheArb_io_mem_resp_bits_replay;
	wire dcacheArb_io_mem_resp_bits_has_data;
	wire [31:0] dcacheArb_io_mem_resp_bits_data_word_bypass;
	wire [31:0] dcacheArb_io_mem_resp_bits_data_raw;
	wire dcacheArb_io_mem_replay_next;
	wire dcacheArb_io_mem_s2_xcpt_ma_ld;
	wire dcacheArb_io_mem_s2_xcpt_ma_st;
	wire dcacheArb_io_mem_s2_xcpt_pf_ld;
	wire dcacheArb_io_mem_s2_xcpt_pf_st;
	wire dcacheArb_io_mem_s2_xcpt_ae_ld;
	wire dcacheArb_io_mem_s2_xcpt_ae_st;
	wire dcacheArb_io_mem_ordered;
	wire dcacheArb_io_mem_perf_grant;
	wire ptw_clock;
	wire ptw_reset;
	wire ptw_io_requestor_0_status_debug;
	wire ptw_io_requestor_0_pmp_0_cfg_l;
	wire [1:0] ptw_io_requestor_0_pmp_0_cfg_a;
	wire ptw_io_requestor_0_pmp_0_cfg_x;
	wire ptw_io_requestor_0_pmp_0_cfg_w;
	wire ptw_io_requestor_0_pmp_0_cfg_r;
	wire [29:0] ptw_io_requestor_0_pmp_0_addr;
	wire [31:0] ptw_io_requestor_0_pmp_0_mask;
	wire ptw_io_requestor_0_pmp_1_cfg_l;
	wire [1:0] ptw_io_requestor_0_pmp_1_cfg_a;
	wire ptw_io_requestor_0_pmp_1_cfg_x;
	wire ptw_io_requestor_0_pmp_1_cfg_w;
	wire ptw_io_requestor_0_pmp_1_cfg_r;
	wire [29:0] ptw_io_requestor_0_pmp_1_addr;
	wire [31:0] ptw_io_requestor_0_pmp_1_mask;
	wire ptw_io_requestor_0_pmp_2_cfg_l;
	wire [1:0] ptw_io_requestor_0_pmp_2_cfg_a;
	wire ptw_io_requestor_0_pmp_2_cfg_x;
	wire ptw_io_requestor_0_pmp_2_cfg_w;
	wire ptw_io_requestor_0_pmp_2_cfg_r;
	wire [29:0] ptw_io_requestor_0_pmp_2_addr;
	wire [31:0] ptw_io_requestor_0_pmp_2_mask;
	wire ptw_io_requestor_0_pmp_3_cfg_l;
	wire [1:0] ptw_io_requestor_0_pmp_3_cfg_a;
	wire ptw_io_requestor_0_pmp_3_cfg_x;
	wire ptw_io_requestor_0_pmp_3_cfg_w;
	wire ptw_io_requestor_0_pmp_3_cfg_r;
	wire [29:0] ptw_io_requestor_0_pmp_3_addr;
	wire [31:0] ptw_io_requestor_0_pmp_3_mask;
	wire ptw_io_requestor_0_pmp_4_cfg_l;
	wire [1:0] ptw_io_requestor_0_pmp_4_cfg_a;
	wire ptw_io_requestor_0_pmp_4_cfg_x;
	wire ptw_io_requestor_0_pmp_4_cfg_w;
	wire ptw_io_requestor_0_pmp_4_cfg_r;
	wire [29:0] ptw_io_requestor_0_pmp_4_addr;
	wire [31:0] ptw_io_requestor_0_pmp_4_mask;
	wire ptw_io_requestor_0_pmp_5_cfg_l;
	wire [1:0] ptw_io_requestor_0_pmp_5_cfg_a;
	wire ptw_io_requestor_0_pmp_5_cfg_x;
	wire ptw_io_requestor_0_pmp_5_cfg_w;
	wire ptw_io_requestor_0_pmp_5_cfg_r;
	wire [29:0] ptw_io_requestor_0_pmp_5_addr;
	wire [31:0] ptw_io_requestor_0_pmp_5_mask;
	wire ptw_io_requestor_0_pmp_6_cfg_l;
	wire [1:0] ptw_io_requestor_0_pmp_6_cfg_a;
	wire ptw_io_requestor_0_pmp_6_cfg_x;
	wire ptw_io_requestor_0_pmp_6_cfg_w;
	wire ptw_io_requestor_0_pmp_6_cfg_r;
	wire [29:0] ptw_io_requestor_0_pmp_6_addr;
	wire [31:0] ptw_io_requestor_0_pmp_6_mask;
	wire ptw_io_requestor_0_pmp_7_cfg_l;
	wire [1:0] ptw_io_requestor_0_pmp_7_cfg_a;
	wire ptw_io_requestor_0_pmp_7_cfg_x;
	wire ptw_io_requestor_0_pmp_7_cfg_w;
	wire ptw_io_requestor_0_pmp_7_cfg_r;
	wire [29:0] ptw_io_requestor_0_pmp_7_addr;
	wire [31:0] ptw_io_requestor_0_pmp_7_mask;
	wire ptw_io_requestor_1_status_debug;
	wire ptw_io_requestor_1_pmp_0_cfg_l;
	wire [1:0] ptw_io_requestor_1_pmp_0_cfg_a;
	wire ptw_io_requestor_1_pmp_0_cfg_x;
	wire ptw_io_requestor_1_pmp_0_cfg_w;
	wire ptw_io_requestor_1_pmp_0_cfg_r;
	wire [29:0] ptw_io_requestor_1_pmp_0_addr;
	wire [31:0] ptw_io_requestor_1_pmp_0_mask;
	wire ptw_io_requestor_1_pmp_1_cfg_l;
	wire [1:0] ptw_io_requestor_1_pmp_1_cfg_a;
	wire ptw_io_requestor_1_pmp_1_cfg_x;
	wire ptw_io_requestor_1_pmp_1_cfg_w;
	wire ptw_io_requestor_1_pmp_1_cfg_r;
	wire [29:0] ptw_io_requestor_1_pmp_1_addr;
	wire [31:0] ptw_io_requestor_1_pmp_1_mask;
	wire ptw_io_requestor_1_pmp_2_cfg_l;
	wire [1:0] ptw_io_requestor_1_pmp_2_cfg_a;
	wire ptw_io_requestor_1_pmp_2_cfg_x;
	wire ptw_io_requestor_1_pmp_2_cfg_w;
	wire ptw_io_requestor_1_pmp_2_cfg_r;
	wire [29:0] ptw_io_requestor_1_pmp_2_addr;
	wire [31:0] ptw_io_requestor_1_pmp_2_mask;
	wire ptw_io_requestor_1_pmp_3_cfg_l;
	wire [1:0] ptw_io_requestor_1_pmp_3_cfg_a;
	wire ptw_io_requestor_1_pmp_3_cfg_x;
	wire ptw_io_requestor_1_pmp_3_cfg_w;
	wire ptw_io_requestor_1_pmp_3_cfg_r;
	wire [29:0] ptw_io_requestor_1_pmp_3_addr;
	wire [31:0] ptw_io_requestor_1_pmp_3_mask;
	wire ptw_io_requestor_1_pmp_4_cfg_l;
	wire [1:0] ptw_io_requestor_1_pmp_4_cfg_a;
	wire ptw_io_requestor_1_pmp_4_cfg_x;
	wire ptw_io_requestor_1_pmp_4_cfg_w;
	wire ptw_io_requestor_1_pmp_4_cfg_r;
	wire [29:0] ptw_io_requestor_1_pmp_4_addr;
	wire [31:0] ptw_io_requestor_1_pmp_4_mask;
	wire ptw_io_requestor_1_pmp_5_cfg_l;
	wire [1:0] ptw_io_requestor_1_pmp_5_cfg_a;
	wire ptw_io_requestor_1_pmp_5_cfg_x;
	wire ptw_io_requestor_1_pmp_5_cfg_w;
	wire ptw_io_requestor_1_pmp_5_cfg_r;
	wire [29:0] ptw_io_requestor_1_pmp_5_addr;
	wire [31:0] ptw_io_requestor_1_pmp_5_mask;
	wire ptw_io_requestor_1_pmp_6_cfg_l;
	wire [1:0] ptw_io_requestor_1_pmp_6_cfg_a;
	wire ptw_io_requestor_1_pmp_6_cfg_x;
	wire ptw_io_requestor_1_pmp_6_cfg_w;
	wire ptw_io_requestor_1_pmp_6_cfg_r;
	wire [29:0] ptw_io_requestor_1_pmp_6_addr;
	wire [31:0] ptw_io_requestor_1_pmp_6_mask;
	wire ptw_io_requestor_1_pmp_7_cfg_l;
	wire [1:0] ptw_io_requestor_1_pmp_7_cfg_a;
	wire ptw_io_requestor_1_pmp_7_cfg_x;
	wire ptw_io_requestor_1_pmp_7_cfg_w;
	wire ptw_io_requestor_1_pmp_7_cfg_r;
	wire [29:0] ptw_io_requestor_1_pmp_7_addr;
	wire [31:0] ptw_io_requestor_1_pmp_7_mask;
	wire [31:0] ptw_io_requestor_1_customCSRs_csrs_0_value;
	wire ptw_io_dpath_status_debug;
	wire ptw_io_dpath_pmp_0_cfg_l;
	wire [1:0] ptw_io_dpath_pmp_0_cfg_a;
	wire ptw_io_dpath_pmp_0_cfg_x;
	wire ptw_io_dpath_pmp_0_cfg_w;
	wire ptw_io_dpath_pmp_0_cfg_r;
	wire [29:0] ptw_io_dpath_pmp_0_addr;
	wire [31:0] ptw_io_dpath_pmp_0_mask;
	wire ptw_io_dpath_pmp_1_cfg_l;
	wire [1:0] ptw_io_dpath_pmp_1_cfg_a;
	wire ptw_io_dpath_pmp_1_cfg_x;
	wire ptw_io_dpath_pmp_1_cfg_w;
	wire ptw_io_dpath_pmp_1_cfg_r;
	wire [29:0] ptw_io_dpath_pmp_1_addr;
	wire [31:0] ptw_io_dpath_pmp_1_mask;
	wire ptw_io_dpath_pmp_2_cfg_l;
	wire [1:0] ptw_io_dpath_pmp_2_cfg_a;
	wire ptw_io_dpath_pmp_2_cfg_x;
	wire ptw_io_dpath_pmp_2_cfg_w;
	wire ptw_io_dpath_pmp_2_cfg_r;
	wire [29:0] ptw_io_dpath_pmp_2_addr;
	wire [31:0] ptw_io_dpath_pmp_2_mask;
	wire ptw_io_dpath_pmp_3_cfg_l;
	wire [1:0] ptw_io_dpath_pmp_3_cfg_a;
	wire ptw_io_dpath_pmp_3_cfg_x;
	wire ptw_io_dpath_pmp_3_cfg_w;
	wire ptw_io_dpath_pmp_3_cfg_r;
	wire [29:0] ptw_io_dpath_pmp_3_addr;
	wire [31:0] ptw_io_dpath_pmp_3_mask;
	wire ptw_io_dpath_pmp_4_cfg_l;
	wire [1:0] ptw_io_dpath_pmp_4_cfg_a;
	wire ptw_io_dpath_pmp_4_cfg_x;
	wire ptw_io_dpath_pmp_4_cfg_w;
	wire ptw_io_dpath_pmp_4_cfg_r;
	wire [29:0] ptw_io_dpath_pmp_4_addr;
	wire [31:0] ptw_io_dpath_pmp_4_mask;
	wire ptw_io_dpath_pmp_5_cfg_l;
	wire [1:0] ptw_io_dpath_pmp_5_cfg_a;
	wire ptw_io_dpath_pmp_5_cfg_x;
	wire ptw_io_dpath_pmp_5_cfg_w;
	wire ptw_io_dpath_pmp_5_cfg_r;
	wire [29:0] ptw_io_dpath_pmp_5_addr;
	wire [31:0] ptw_io_dpath_pmp_5_mask;
	wire ptw_io_dpath_pmp_6_cfg_l;
	wire [1:0] ptw_io_dpath_pmp_6_cfg_a;
	wire ptw_io_dpath_pmp_6_cfg_x;
	wire ptw_io_dpath_pmp_6_cfg_w;
	wire ptw_io_dpath_pmp_6_cfg_r;
	wire [29:0] ptw_io_dpath_pmp_6_addr;
	wire [31:0] ptw_io_dpath_pmp_6_mask;
	wire ptw_io_dpath_pmp_7_cfg_l;
	wire [1:0] ptw_io_dpath_pmp_7_cfg_a;
	wire ptw_io_dpath_pmp_7_cfg_x;
	wire ptw_io_dpath_pmp_7_cfg_w;
	wire ptw_io_dpath_pmp_7_cfg_r;
	wire [29:0] ptw_io_dpath_pmp_7_addr;
	wire [31:0] ptw_io_dpath_pmp_7_mask;
	wire ptw_io_dpath_perf_l2hit;
	wire ptw_io_dpath_perf_pte_miss;
	wire ptw_io_dpath_perf_pte_hit;
	wire [31:0] ptw_io_dpath_customCSRs_csrs_0_value;
	wire core_clock;
	wire core_reset;
	wire core_io_hartid;
	wire core_io_interrupts_debug;
	wire core_io_interrupts_mtip;
	wire core_io_interrupts_msip;
	wire core_io_interrupts_meip;
	wire core_io_imem_might_request;
	wire core_io_imem_req_valid;
	wire [31:0] core_io_imem_req_bits_pc;
	wire core_io_imem_req_bits_speculative;
	wire core_io_imem_resp_ready;
	wire core_io_imem_resp_valid;
	wire [31:0] core_io_imem_resp_bits_pc;
	wire [31:0] core_io_imem_resp_bits_data;
	wire core_io_imem_resp_bits_xcpt_ae_inst;
	wire core_io_imem_resp_bits_replay;
	wire core_io_imem_btb_update_valid;
	wire core_io_imem_bht_update_valid;
	wire core_io_imem_flush_icache;
	wire core_io_dmem_req_ready;
	wire core_io_dmem_req_valid;
	wire [31:0] core_io_dmem_req_bits_addr;
	wire [6:0] core_io_dmem_req_bits_tag;
	wire [4:0] core_io_dmem_req_bits_cmd;
	wire [1:0] core_io_dmem_req_bits_size;
	wire core_io_dmem_req_bits_signed;
	wire core_io_dmem_req_bits_dv;
	wire core_io_dmem_s1_kill;
	wire [31:0] core_io_dmem_s1_data_data;
	wire core_io_dmem_s2_nack;
	wire core_io_dmem_resp_valid;
	wire [6:0] core_io_dmem_resp_bits_tag;
	wire [31:0] core_io_dmem_resp_bits_data;
	wire core_io_dmem_resp_bits_replay;
	wire core_io_dmem_resp_bits_has_data;
	wire [31:0] core_io_dmem_resp_bits_data_word_bypass;
	wire core_io_dmem_replay_next;
	wire core_io_dmem_s2_xcpt_ma_ld;
	wire core_io_dmem_s2_xcpt_ma_st;
	wire core_io_dmem_s2_xcpt_pf_ld;
	wire core_io_dmem_s2_xcpt_pf_st;
	wire core_io_dmem_s2_xcpt_ae_ld;
	wire core_io_dmem_s2_xcpt_ae_st;
	wire core_io_dmem_ordered;
	wire core_io_dmem_perf_grant;
	wire core_io_ptw_status_debug;
	wire core_io_ptw_pmp_0_cfg_l;
	wire [1:0] core_io_ptw_pmp_0_cfg_a;
	wire core_io_ptw_pmp_0_cfg_x;
	wire core_io_ptw_pmp_0_cfg_w;
	wire core_io_ptw_pmp_0_cfg_r;
	wire [29:0] core_io_ptw_pmp_0_addr;
	wire [31:0] core_io_ptw_pmp_0_mask;
	wire core_io_ptw_pmp_1_cfg_l;
	wire [1:0] core_io_ptw_pmp_1_cfg_a;
	wire core_io_ptw_pmp_1_cfg_x;
	wire core_io_ptw_pmp_1_cfg_w;
	wire core_io_ptw_pmp_1_cfg_r;
	wire [29:0] core_io_ptw_pmp_1_addr;
	wire [31:0] core_io_ptw_pmp_1_mask;
	wire core_io_ptw_pmp_2_cfg_l;
	wire [1:0] core_io_ptw_pmp_2_cfg_a;
	wire core_io_ptw_pmp_2_cfg_x;
	wire core_io_ptw_pmp_2_cfg_w;
	wire core_io_ptw_pmp_2_cfg_r;
	wire [29:0] core_io_ptw_pmp_2_addr;
	wire [31:0] core_io_ptw_pmp_2_mask;
	wire core_io_ptw_pmp_3_cfg_l;
	wire [1:0] core_io_ptw_pmp_3_cfg_a;
	wire core_io_ptw_pmp_3_cfg_x;
	wire core_io_ptw_pmp_3_cfg_w;
	wire core_io_ptw_pmp_3_cfg_r;
	wire [29:0] core_io_ptw_pmp_3_addr;
	wire [31:0] core_io_ptw_pmp_3_mask;
	wire core_io_ptw_pmp_4_cfg_l;
	wire [1:0] core_io_ptw_pmp_4_cfg_a;
	wire core_io_ptw_pmp_4_cfg_x;
	wire core_io_ptw_pmp_4_cfg_w;
	wire core_io_ptw_pmp_4_cfg_r;
	wire [29:0] core_io_ptw_pmp_4_addr;
	wire [31:0] core_io_ptw_pmp_4_mask;
	wire core_io_ptw_pmp_5_cfg_l;
	wire [1:0] core_io_ptw_pmp_5_cfg_a;
	wire core_io_ptw_pmp_5_cfg_x;
	wire core_io_ptw_pmp_5_cfg_w;
	wire core_io_ptw_pmp_5_cfg_r;
	wire [29:0] core_io_ptw_pmp_5_addr;
	wire [31:0] core_io_ptw_pmp_5_mask;
	wire core_io_ptw_pmp_6_cfg_l;
	wire [1:0] core_io_ptw_pmp_6_cfg_a;
	wire core_io_ptw_pmp_6_cfg_x;
	wire core_io_ptw_pmp_6_cfg_w;
	wire core_io_ptw_pmp_6_cfg_r;
	wire [29:0] core_io_ptw_pmp_6_addr;
	wire [31:0] core_io_ptw_pmp_6_mask;
	wire core_io_ptw_pmp_7_cfg_l;
	wire [1:0] core_io_ptw_pmp_7_cfg_a;
	wire core_io_ptw_pmp_7_cfg_x;
	wire core_io_ptw_pmp_7_cfg_w;
	wire core_io_ptw_pmp_7_cfg_r;
	wire [29:0] core_io_ptw_pmp_7_addr;
	wire [31:0] core_io_ptw_pmp_7_mask;
	wire [31:0] core_io_ptw_customCSRs_csrs_0_value;
	wire core_io_wfi;
	reg bundleOut_0_0_REG;
	TLXbar_6 tlMasterXbar(
		.clock(tlMasterXbar_clock),
		.reset(tlMasterXbar_reset),
		.auto_in_1_a_ready(tlMasterXbar_auto_in_1_a_ready),
		.auto_in_1_a_valid(tlMasterXbar_auto_in_1_a_valid),
		.auto_in_1_a_bits_address(tlMasterXbar_auto_in_1_a_bits_address),
		.auto_in_1_d_valid(tlMasterXbar_auto_in_1_d_valid),
		.auto_in_1_d_bits_opcode(tlMasterXbar_auto_in_1_d_bits_opcode),
		.auto_in_1_d_bits_size(tlMasterXbar_auto_in_1_d_bits_size),
		.auto_in_1_d_bits_data(tlMasterXbar_auto_in_1_d_bits_data),
		.auto_in_1_d_bits_corrupt(tlMasterXbar_auto_in_1_d_bits_corrupt),
		.auto_in_0_a_ready(tlMasterXbar_auto_in_0_a_ready),
		.auto_in_0_a_valid(tlMasterXbar_auto_in_0_a_valid),
		.auto_in_0_a_bits_opcode(tlMasterXbar_auto_in_0_a_bits_opcode),
		.auto_in_0_a_bits_param(tlMasterXbar_auto_in_0_a_bits_param),
		.auto_in_0_a_bits_size(tlMasterXbar_auto_in_0_a_bits_size),
		.auto_in_0_a_bits_address(tlMasterXbar_auto_in_0_a_bits_address),
		.auto_in_0_a_bits_mask(tlMasterXbar_auto_in_0_a_bits_mask),
		.auto_in_0_a_bits_data(tlMasterXbar_auto_in_0_a_bits_data),
		.auto_in_0_d_ready(tlMasterXbar_auto_in_0_d_ready),
		.auto_in_0_d_valid(tlMasterXbar_auto_in_0_d_valid),
		.auto_in_0_d_bits_opcode(tlMasterXbar_auto_in_0_d_bits_opcode),
		.auto_in_0_d_bits_size(tlMasterXbar_auto_in_0_d_bits_size),
		.auto_in_0_d_bits_denied(tlMasterXbar_auto_in_0_d_bits_denied),
		.auto_in_0_d_bits_data(tlMasterXbar_auto_in_0_d_bits_data),
		.auto_out_a_ready(tlMasterXbar_auto_out_a_ready),
		.auto_out_a_valid(tlMasterXbar_auto_out_a_valid),
		.auto_out_a_bits_opcode(tlMasterXbar_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(tlMasterXbar_auto_out_a_bits_param),
		.auto_out_a_bits_size(tlMasterXbar_auto_out_a_bits_size),
		.auto_out_a_bits_source(tlMasterXbar_auto_out_a_bits_source),
		.auto_out_a_bits_address(tlMasterXbar_auto_out_a_bits_address),
		.auto_out_a_bits_mask(tlMasterXbar_auto_out_a_bits_mask),
		.auto_out_a_bits_data(tlMasterXbar_auto_out_a_bits_data),
		.auto_out_d_ready(tlMasterXbar_auto_out_d_ready),
		.auto_out_d_valid(tlMasterXbar_auto_out_d_valid),
		.auto_out_d_bits_opcode(tlMasterXbar_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(tlMasterXbar_auto_out_d_bits_param),
		.auto_out_d_bits_size(tlMasterXbar_auto_out_d_bits_size),
		.auto_out_d_bits_source(tlMasterXbar_auto_out_d_bits_source),
		.auto_out_d_bits_sink(tlMasterXbar_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(tlMasterXbar_auto_out_d_bits_denied),
		.auto_out_d_bits_data(tlMasterXbar_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(tlMasterXbar_auto_out_d_bits_corrupt)
	);
	TLXbar_7 tlSlaveXbar(
		.auto_in_a_ready(tlSlaveXbar_auto_in_a_ready),
		.auto_in_a_valid(tlSlaveXbar_auto_in_a_valid),
		.auto_in_a_bits_opcode(tlSlaveXbar_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(tlSlaveXbar_auto_in_a_bits_param),
		.auto_in_a_bits_size(tlSlaveXbar_auto_in_a_bits_size),
		.auto_in_a_bits_source(tlSlaveXbar_auto_in_a_bits_source),
		.auto_in_a_bits_address(tlSlaveXbar_auto_in_a_bits_address),
		.auto_in_a_bits_mask(tlSlaveXbar_auto_in_a_bits_mask),
		.auto_in_a_bits_data(tlSlaveXbar_auto_in_a_bits_data),
		.auto_in_d_ready(tlSlaveXbar_auto_in_d_ready),
		.auto_in_d_valid(tlSlaveXbar_auto_in_d_valid),
		.auto_in_d_bits_opcode(tlSlaveXbar_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(tlSlaveXbar_auto_in_d_bits_size),
		.auto_in_d_bits_source(tlSlaveXbar_auto_in_d_bits_source),
		.auto_in_d_bits_data(tlSlaveXbar_auto_in_d_bits_data),
		.auto_out_a_ready(tlSlaveXbar_auto_out_a_ready),
		.auto_out_a_valid(tlSlaveXbar_auto_out_a_valid),
		.auto_out_a_bits_opcode(tlSlaveXbar_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(tlSlaveXbar_auto_out_a_bits_param),
		.auto_out_a_bits_size(tlSlaveXbar_auto_out_a_bits_size),
		.auto_out_a_bits_source(tlSlaveXbar_auto_out_a_bits_source),
		.auto_out_a_bits_address(tlSlaveXbar_auto_out_a_bits_address),
		.auto_out_a_bits_mask(tlSlaveXbar_auto_out_a_bits_mask),
		.auto_out_a_bits_data(tlSlaveXbar_auto_out_a_bits_data),
		.auto_out_d_ready(tlSlaveXbar_auto_out_d_ready),
		.auto_out_d_valid(tlSlaveXbar_auto_out_d_valid),
		.auto_out_d_bits_opcode(tlSlaveXbar_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(tlSlaveXbar_auto_out_d_bits_size),
		.auto_out_d_bits_source(tlSlaveXbar_auto_out_d_bits_source),
		.auto_out_d_bits_data(tlSlaveXbar_auto_out_d_bits_data)
	);
	IntXbar_1 intXbar(
		.auto_int_in_2_0(intXbar_auto_int_in_2_0),
		.auto_int_in_1_0(intXbar_auto_int_in_1_0),
		.auto_int_in_1_1(intXbar_auto_int_in_1_1),
		.auto_int_in_0_0(intXbar_auto_int_in_0_0),
		.auto_int_out_0(intXbar_auto_int_out_0),
		.auto_int_out_1(intXbar_auto_int_out_1),
		.auto_int_out_2(intXbar_auto_int_out_2),
		.auto_int_out_3(intXbar_auto_int_out_3)
	);
	BundleBridgeNexus_4 broadcast(
		.auto_in(broadcast_auto_in),
		.auto_out_0(broadcast_auto_out_0)
	);
	DCache dcache(
		.clock(dcache_clock),
		.reset(dcache_reset),
		.auto_out_a_ready(dcache_auto_out_a_ready),
		.auto_out_a_valid(dcache_auto_out_a_valid),
		.auto_out_a_bits_opcode(dcache_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(dcache_auto_out_a_bits_param),
		.auto_out_a_bits_size(dcache_auto_out_a_bits_size),
		.auto_out_a_bits_address(dcache_auto_out_a_bits_address),
		.auto_out_a_bits_mask(dcache_auto_out_a_bits_mask),
		.auto_out_a_bits_data(dcache_auto_out_a_bits_data),
		.auto_out_d_ready(dcache_auto_out_d_ready),
		.auto_out_d_valid(dcache_auto_out_d_valid),
		.auto_out_d_bits_opcode(dcache_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(dcache_auto_out_d_bits_size),
		.auto_out_d_bits_denied(dcache_auto_out_d_bits_denied),
		.auto_out_d_bits_data(dcache_auto_out_d_bits_data),
		.io_cpu_req_ready(dcache_io_cpu_req_ready),
		.io_cpu_req_valid(dcache_io_cpu_req_valid),
		.io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr),
		.io_cpu_req_bits_tag(dcache_io_cpu_req_bits_tag),
		.io_cpu_req_bits_cmd(dcache_io_cpu_req_bits_cmd),
		.io_cpu_req_bits_size(dcache_io_cpu_req_bits_size),
		.io_cpu_req_bits_signed(dcache_io_cpu_req_bits_signed),
		.io_cpu_req_bits_dprv(dcache_io_cpu_req_bits_dprv),
		.io_cpu_req_bits_no_xcpt(dcache_io_cpu_req_bits_no_xcpt),
		.io_cpu_s1_kill(dcache_io_cpu_s1_kill),
		.io_cpu_s1_data_data(dcache_io_cpu_s1_data_data),
		.io_cpu_s1_data_mask(dcache_io_cpu_s1_data_mask),
		.io_cpu_s2_nack(dcache_io_cpu_s2_nack),
		.io_cpu_resp_valid(dcache_io_cpu_resp_valid),
		.io_cpu_resp_bits_addr(dcache_io_cpu_resp_bits_addr),
		.io_cpu_resp_bits_tag(dcache_io_cpu_resp_bits_tag),
		.io_cpu_resp_bits_cmd(dcache_io_cpu_resp_bits_cmd),
		.io_cpu_resp_bits_size(dcache_io_cpu_resp_bits_size),
		.io_cpu_resp_bits_signed(dcache_io_cpu_resp_bits_signed),
		.io_cpu_resp_bits_dprv(dcache_io_cpu_resp_bits_dprv),
		.io_cpu_resp_bits_dv(dcache_io_cpu_resp_bits_dv),
		.io_cpu_resp_bits_data(dcache_io_cpu_resp_bits_data),
		.io_cpu_resp_bits_mask(dcache_io_cpu_resp_bits_mask),
		.io_cpu_resp_bits_replay(dcache_io_cpu_resp_bits_replay),
		.io_cpu_resp_bits_has_data(dcache_io_cpu_resp_bits_has_data),
		.io_cpu_resp_bits_data_word_bypass(dcache_io_cpu_resp_bits_data_word_bypass),
		.io_cpu_resp_bits_data_raw(dcache_io_cpu_resp_bits_data_raw),
		.io_cpu_resp_bits_store_data(dcache_io_cpu_resp_bits_store_data),
		.io_cpu_replay_next(dcache_io_cpu_replay_next),
		.io_cpu_s2_xcpt_ma_ld(dcache_io_cpu_s2_xcpt_ma_ld),
		.io_cpu_s2_xcpt_ma_st(dcache_io_cpu_s2_xcpt_ma_st),
		.io_cpu_s2_xcpt_pf_ld(dcache_io_cpu_s2_xcpt_pf_ld),
		.io_cpu_s2_xcpt_pf_st(dcache_io_cpu_s2_xcpt_pf_st),
		.io_cpu_s2_xcpt_gf_ld(dcache_io_cpu_s2_xcpt_gf_ld),
		.io_cpu_s2_xcpt_gf_st(dcache_io_cpu_s2_xcpt_gf_st),
		.io_cpu_s2_xcpt_ae_ld(dcache_io_cpu_s2_xcpt_ae_ld),
		.io_cpu_s2_xcpt_ae_st(dcache_io_cpu_s2_xcpt_ae_st),
		.io_cpu_ordered(dcache_io_cpu_ordered),
		.io_cpu_perf_grant(dcache_io_cpu_perf_grant),
		.io_ptw_status_debug(dcache_io_ptw_status_debug),
		.io_ptw_pmp_0_cfg_l(dcache_io_ptw_pmp_0_cfg_l),
		.io_ptw_pmp_0_cfg_a(dcache_io_ptw_pmp_0_cfg_a),
		.io_ptw_pmp_0_cfg_x(dcache_io_ptw_pmp_0_cfg_x),
		.io_ptw_pmp_0_cfg_w(dcache_io_ptw_pmp_0_cfg_w),
		.io_ptw_pmp_0_cfg_r(dcache_io_ptw_pmp_0_cfg_r),
		.io_ptw_pmp_0_addr(dcache_io_ptw_pmp_0_addr),
		.io_ptw_pmp_0_mask(dcache_io_ptw_pmp_0_mask),
		.io_ptw_pmp_1_cfg_l(dcache_io_ptw_pmp_1_cfg_l),
		.io_ptw_pmp_1_cfg_a(dcache_io_ptw_pmp_1_cfg_a),
		.io_ptw_pmp_1_cfg_x(dcache_io_ptw_pmp_1_cfg_x),
		.io_ptw_pmp_1_cfg_w(dcache_io_ptw_pmp_1_cfg_w),
		.io_ptw_pmp_1_cfg_r(dcache_io_ptw_pmp_1_cfg_r),
		.io_ptw_pmp_1_addr(dcache_io_ptw_pmp_1_addr),
		.io_ptw_pmp_1_mask(dcache_io_ptw_pmp_1_mask),
		.io_ptw_pmp_2_cfg_l(dcache_io_ptw_pmp_2_cfg_l),
		.io_ptw_pmp_2_cfg_a(dcache_io_ptw_pmp_2_cfg_a),
		.io_ptw_pmp_2_cfg_x(dcache_io_ptw_pmp_2_cfg_x),
		.io_ptw_pmp_2_cfg_w(dcache_io_ptw_pmp_2_cfg_w),
		.io_ptw_pmp_2_cfg_r(dcache_io_ptw_pmp_2_cfg_r),
		.io_ptw_pmp_2_addr(dcache_io_ptw_pmp_2_addr),
		.io_ptw_pmp_2_mask(dcache_io_ptw_pmp_2_mask),
		.io_ptw_pmp_3_cfg_l(dcache_io_ptw_pmp_3_cfg_l),
		.io_ptw_pmp_3_cfg_a(dcache_io_ptw_pmp_3_cfg_a),
		.io_ptw_pmp_3_cfg_x(dcache_io_ptw_pmp_3_cfg_x),
		.io_ptw_pmp_3_cfg_w(dcache_io_ptw_pmp_3_cfg_w),
		.io_ptw_pmp_3_cfg_r(dcache_io_ptw_pmp_3_cfg_r),
		.io_ptw_pmp_3_addr(dcache_io_ptw_pmp_3_addr),
		.io_ptw_pmp_3_mask(dcache_io_ptw_pmp_3_mask),
		.io_ptw_pmp_4_cfg_l(dcache_io_ptw_pmp_4_cfg_l),
		.io_ptw_pmp_4_cfg_a(dcache_io_ptw_pmp_4_cfg_a),
		.io_ptw_pmp_4_cfg_x(dcache_io_ptw_pmp_4_cfg_x),
		.io_ptw_pmp_4_cfg_w(dcache_io_ptw_pmp_4_cfg_w),
		.io_ptw_pmp_4_cfg_r(dcache_io_ptw_pmp_4_cfg_r),
		.io_ptw_pmp_4_addr(dcache_io_ptw_pmp_4_addr),
		.io_ptw_pmp_4_mask(dcache_io_ptw_pmp_4_mask),
		.io_ptw_pmp_5_cfg_l(dcache_io_ptw_pmp_5_cfg_l),
		.io_ptw_pmp_5_cfg_a(dcache_io_ptw_pmp_5_cfg_a),
		.io_ptw_pmp_5_cfg_x(dcache_io_ptw_pmp_5_cfg_x),
		.io_ptw_pmp_5_cfg_w(dcache_io_ptw_pmp_5_cfg_w),
		.io_ptw_pmp_5_cfg_r(dcache_io_ptw_pmp_5_cfg_r),
		.io_ptw_pmp_5_addr(dcache_io_ptw_pmp_5_addr),
		.io_ptw_pmp_5_mask(dcache_io_ptw_pmp_5_mask),
		.io_ptw_pmp_6_cfg_l(dcache_io_ptw_pmp_6_cfg_l),
		.io_ptw_pmp_6_cfg_a(dcache_io_ptw_pmp_6_cfg_a),
		.io_ptw_pmp_6_cfg_x(dcache_io_ptw_pmp_6_cfg_x),
		.io_ptw_pmp_6_cfg_w(dcache_io_ptw_pmp_6_cfg_w),
		.io_ptw_pmp_6_cfg_r(dcache_io_ptw_pmp_6_cfg_r),
		.io_ptw_pmp_6_addr(dcache_io_ptw_pmp_6_addr),
		.io_ptw_pmp_6_mask(dcache_io_ptw_pmp_6_mask),
		.io_ptw_pmp_7_cfg_l(dcache_io_ptw_pmp_7_cfg_l),
		.io_ptw_pmp_7_cfg_a(dcache_io_ptw_pmp_7_cfg_a),
		.io_ptw_pmp_7_cfg_x(dcache_io_ptw_pmp_7_cfg_x),
		.io_ptw_pmp_7_cfg_w(dcache_io_ptw_pmp_7_cfg_w),
		.io_ptw_pmp_7_cfg_r(dcache_io_ptw_pmp_7_cfg_r),
		.io_ptw_pmp_7_addr(dcache_io_ptw_pmp_7_addr),
		.io_ptw_pmp_7_mask(dcache_io_ptw_pmp_7_mask)
	);
	Frontend frontend(
		.clock(frontend_clock),
		.reset(frontend_reset),
		.auto_icache_master_out_a_ready(frontend_auto_icache_master_out_a_ready),
		.auto_icache_master_out_a_valid(frontend_auto_icache_master_out_a_valid),
		.auto_icache_master_out_a_bits_address(frontend_auto_icache_master_out_a_bits_address),
		.auto_icache_master_out_d_valid(frontend_auto_icache_master_out_d_valid),
		.auto_icache_master_out_d_bits_opcode(frontend_auto_icache_master_out_d_bits_opcode),
		.auto_icache_master_out_d_bits_size(frontend_auto_icache_master_out_d_bits_size),
		.auto_icache_master_out_d_bits_data(frontend_auto_icache_master_out_d_bits_data),
		.auto_icache_master_out_d_bits_corrupt(frontend_auto_icache_master_out_d_bits_corrupt),
		.io_cpu_might_request(frontend_io_cpu_might_request),
		.io_cpu_req_valid(frontend_io_cpu_req_valid),
		.io_cpu_req_bits_pc(frontend_io_cpu_req_bits_pc),
		.io_cpu_req_bits_speculative(frontend_io_cpu_req_bits_speculative),
		.io_cpu_resp_ready(frontend_io_cpu_resp_ready),
		.io_cpu_resp_valid(frontend_io_cpu_resp_valid),
		.io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),
		.io_cpu_resp_bits_data(frontend_io_cpu_resp_bits_data),
		.io_cpu_resp_bits_xcpt_ae_inst(frontend_io_cpu_resp_bits_xcpt_ae_inst),
		.io_cpu_resp_bits_replay(frontend_io_cpu_resp_bits_replay),
		.io_cpu_btb_update_valid(frontend_io_cpu_btb_update_valid),
		.io_cpu_bht_update_valid(frontend_io_cpu_bht_update_valid),
		.io_cpu_flush_icache(frontend_io_cpu_flush_icache),
		.io_cpu_npc(frontend_io_cpu_npc),
		.io_ptw_status_debug(frontend_io_ptw_status_debug),
		.io_ptw_pmp_0_cfg_l(frontend_io_ptw_pmp_0_cfg_l),
		.io_ptw_pmp_0_cfg_a(frontend_io_ptw_pmp_0_cfg_a),
		.io_ptw_pmp_0_cfg_x(frontend_io_ptw_pmp_0_cfg_x),
		.io_ptw_pmp_0_cfg_w(frontend_io_ptw_pmp_0_cfg_w),
		.io_ptw_pmp_0_cfg_r(frontend_io_ptw_pmp_0_cfg_r),
		.io_ptw_pmp_0_addr(frontend_io_ptw_pmp_0_addr),
		.io_ptw_pmp_0_mask(frontend_io_ptw_pmp_0_mask),
		.io_ptw_pmp_1_cfg_l(frontend_io_ptw_pmp_1_cfg_l),
		.io_ptw_pmp_1_cfg_a(frontend_io_ptw_pmp_1_cfg_a),
		.io_ptw_pmp_1_cfg_x(frontend_io_ptw_pmp_1_cfg_x),
		.io_ptw_pmp_1_cfg_w(frontend_io_ptw_pmp_1_cfg_w),
		.io_ptw_pmp_1_cfg_r(frontend_io_ptw_pmp_1_cfg_r),
		.io_ptw_pmp_1_addr(frontend_io_ptw_pmp_1_addr),
		.io_ptw_pmp_1_mask(frontend_io_ptw_pmp_1_mask),
		.io_ptw_pmp_2_cfg_l(frontend_io_ptw_pmp_2_cfg_l),
		.io_ptw_pmp_2_cfg_a(frontend_io_ptw_pmp_2_cfg_a),
		.io_ptw_pmp_2_cfg_x(frontend_io_ptw_pmp_2_cfg_x),
		.io_ptw_pmp_2_cfg_w(frontend_io_ptw_pmp_2_cfg_w),
		.io_ptw_pmp_2_cfg_r(frontend_io_ptw_pmp_2_cfg_r),
		.io_ptw_pmp_2_addr(frontend_io_ptw_pmp_2_addr),
		.io_ptw_pmp_2_mask(frontend_io_ptw_pmp_2_mask),
		.io_ptw_pmp_3_cfg_l(frontend_io_ptw_pmp_3_cfg_l),
		.io_ptw_pmp_3_cfg_a(frontend_io_ptw_pmp_3_cfg_a),
		.io_ptw_pmp_3_cfg_x(frontend_io_ptw_pmp_3_cfg_x),
		.io_ptw_pmp_3_cfg_w(frontend_io_ptw_pmp_3_cfg_w),
		.io_ptw_pmp_3_cfg_r(frontend_io_ptw_pmp_3_cfg_r),
		.io_ptw_pmp_3_addr(frontend_io_ptw_pmp_3_addr),
		.io_ptw_pmp_3_mask(frontend_io_ptw_pmp_3_mask),
		.io_ptw_pmp_4_cfg_l(frontend_io_ptw_pmp_4_cfg_l),
		.io_ptw_pmp_4_cfg_a(frontend_io_ptw_pmp_4_cfg_a),
		.io_ptw_pmp_4_cfg_x(frontend_io_ptw_pmp_4_cfg_x),
		.io_ptw_pmp_4_cfg_w(frontend_io_ptw_pmp_4_cfg_w),
		.io_ptw_pmp_4_cfg_r(frontend_io_ptw_pmp_4_cfg_r),
		.io_ptw_pmp_4_addr(frontend_io_ptw_pmp_4_addr),
		.io_ptw_pmp_4_mask(frontend_io_ptw_pmp_4_mask),
		.io_ptw_pmp_5_cfg_l(frontend_io_ptw_pmp_5_cfg_l),
		.io_ptw_pmp_5_cfg_a(frontend_io_ptw_pmp_5_cfg_a),
		.io_ptw_pmp_5_cfg_x(frontend_io_ptw_pmp_5_cfg_x),
		.io_ptw_pmp_5_cfg_w(frontend_io_ptw_pmp_5_cfg_w),
		.io_ptw_pmp_5_cfg_r(frontend_io_ptw_pmp_5_cfg_r),
		.io_ptw_pmp_5_addr(frontend_io_ptw_pmp_5_addr),
		.io_ptw_pmp_5_mask(frontend_io_ptw_pmp_5_mask),
		.io_ptw_pmp_6_cfg_l(frontend_io_ptw_pmp_6_cfg_l),
		.io_ptw_pmp_6_cfg_a(frontend_io_ptw_pmp_6_cfg_a),
		.io_ptw_pmp_6_cfg_x(frontend_io_ptw_pmp_6_cfg_x),
		.io_ptw_pmp_6_cfg_w(frontend_io_ptw_pmp_6_cfg_w),
		.io_ptw_pmp_6_cfg_r(frontend_io_ptw_pmp_6_cfg_r),
		.io_ptw_pmp_6_addr(frontend_io_ptw_pmp_6_addr),
		.io_ptw_pmp_6_mask(frontend_io_ptw_pmp_6_mask),
		.io_ptw_pmp_7_cfg_l(frontend_io_ptw_pmp_7_cfg_l),
		.io_ptw_pmp_7_cfg_a(frontend_io_ptw_pmp_7_cfg_a),
		.io_ptw_pmp_7_cfg_x(frontend_io_ptw_pmp_7_cfg_x),
		.io_ptw_pmp_7_cfg_w(frontend_io_ptw_pmp_7_cfg_w),
		.io_ptw_pmp_7_cfg_r(frontend_io_ptw_pmp_7_cfg_r),
		.io_ptw_pmp_7_addr(frontend_io_ptw_pmp_7_addr),
		.io_ptw_pmp_7_mask(frontend_io_ptw_pmp_7_mask),
		.io_ptw_customCSRs_csrs_0_value(frontend_io_ptw_customCSRs_csrs_0_value)
	);
	ScratchpadSlavePort dtim_adapter(
		.clock(dtim_adapter_clock),
		.reset(dtim_adapter_reset),
		.auto_in_a_ready(dtim_adapter_auto_in_a_ready),
		.auto_in_a_valid(dtim_adapter_auto_in_a_valid),
		.auto_in_a_bits_opcode(dtim_adapter_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(dtim_adapter_auto_in_a_bits_param),
		.auto_in_a_bits_size(dtim_adapter_auto_in_a_bits_size),
		.auto_in_a_bits_source(dtim_adapter_auto_in_a_bits_source),
		.auto_in_a_bits_address(dtim_adapter_auto_in_a_bits_address),
		.auto_in_a_bits_mask(dtim_adapter_auto_in_a_bits_mask),
		.auto_in_a_bits_data(dtim_adapter_auto_in_a_bits_data),
		.auto_in_d_ready(dtim_adapter_auto_in_d_ready),
		.auto_in_d_valid(dtim_adapter_auto_in_d_valid),
		.auto_in_d_bits_opcode(dtim_adapter_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(dtim_adapter_auto_in_d_bits_size),
		.auto_in_d_bits_source(dtim_adapter_auto_in_d_bits_source),
		.auto_in_d_bits_data(dtim_adapter_auto_in_d_bits_data),
		.io_dmem_req_ready(dtim_adapter_io_dmem_req_ready),
		.io_dmem_req_valid(dtim_adapter_io_dmem_req_valid),
		.io_dmem_req_bits_addr(dtim_adapter_io_dmem_req_bits_addr),
		.io_dmem_req_bits_cmd(dtim_adapter_io_dmem_req_bits_cmd),
		.io_dmem_req_bits_size(dtim_adapter_io_dmem_req_bits_size),
		.io_dmem_s1_kill(dtim_adapter_io_dmem_s1_kill),
		.io_dmem_s1_data_data(dtim_adapter_io_dmem_s1_data_data),
		.io_dmem_s1_data_mask(dtim_adapter_io_dmem_s1_data_mask),
		.io_dmem_s2_nack(dtim_adapter_io_dmem_s2_nack),
		.io_dmem_resp_valid(dtim_adapter_io_dmem_resp_valid),
		.io_dmem_resp_bits_data_raw(dtim_adapter_io_dmem_resp_bits_data_raw)
	);
	TLFragmenter_9 fragmenter_1(
		.clock(fragmenter_1_clock),
		.reset(fragmenter_1_reset),
		.auto_in_a_ready(fragmenter_1_auto_in_a_ready),
		.auto_in_a_valid(fragmenter_1_auto_in_a_valid),
		.auto_in_a_bits_opcode(fragmenter_1_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(fragmenter_1_auto_in_a_bits_param),
		.auto_in_a_bits_size(fragmenter_1_auto_in_a_bits_size),
		.auto_in_a_bits_source(fragmenter_1_auto_in_a_bits_source),
		.auto_in_a_bits_address(fragmenter_1_auto_in_a_bits_address),
		.auto_in_a_bits_mask(fragmenter_1_auto_in_a_bits_mask),
		.auto_in_a_bits_data(fragmenter_1_auto_in_a_bits_data),
		.auto_in_d_ready(fragmenter_1_auto_in_d_ready),
		.auto_in_d_valid(fragmenter_1_auto_in_d_valid),
		.auto_in_d_bits_opcode(fragmenter_1_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(fragmenter_1_auto_in_d_bits_size),
		.auto_in_d_bits_source(fragmenter_1_auto_in_d_bits_source),
		.auto_in_d_bits_data(fragmenter_1_auto_in_d_bits_data),
		.auto_out_a_ready(fragmenter_1_auto_out_a_ready),
		.auto_out_a_valid(fragmenter_1_auto_out_a_valid),
		.auto_out_a_bits_opcode(fragmenter_1_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(fragmenter_1_auto_out_a_bits_param),
		.auto_out_a_bits_size(fragmenter_1_auto_out_a_bits_size),
		.auto_out_a_bits_source(fragmenter_1_auto_out_a_bits_source),
		.auto_out_a_bits_address(fragmenter_1_auto_out_a_bits_address),
		.auto_out_a_bits_mask(fragmenter_1_auto_out_a_bits_mask),
		.auto_out_a_bits_data(fragmenter_1_auto_out_a_bits_data),
		.auto_out_d_ready(fragmenter_1_auto_out_d_ready),
		.auto_out_d_valid(fragmenter_1_auto_out_d_valid),
		.auto_out_d_bits_opcode(fragmenter_1_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(fragmenter_1_auto_out_d_bits_size),
		.auto_out_d_bits_source(fragmenter_1_auto_out_d_bits_source),
		.auto_out_d_bits_data(fragmenter_1_auto_out_d_bits_data)
	);
	HellaCacheArbiter dcacheArb(
		.clock(dcacheArb_clock),
		.io_requestor_0_req_ready(dcacheArb_io_requestor_0_req_ready),
		.io_requestor_0_req_valid(dcacheArb_io_requestor_0_req_valid),
		.io_requestor_0_req_bits_addr(dcacheArb_io_requestor_0_req_bits_addr),
		.io_requestor_0_req_bits_tag(dcacheArb_io_requestor_0_req_bits_tag),
		.io_requestor_0_req_bits_cmd(dcacheArb_io_requestor_0_req_bits_cmd),
		.io_requestor_0_req_bits_size(dcacheArb_io_requestor_0_req_bits_size),
		.io_requestor_0_req_bits_signed(dcacheArb_io_requestor_0_req_bits_signed),
		.io_requestor_0_s1_kill(dcacheArb_io_requestor_0_s1_kill),
		.io_requestor_0_s1_data_data(dcacheArb_io_requestor_0_s1_data_data),
		.io_requestor_0_s2_nack(dcacheArb_io_requestor_0_s2_nack),
		.io_requestor_0_resp_valid(dcacheArb_io_requestor_0_resp_valid),
		.io_requestor_0_resp_bits_tag(dcacheArb_io_requestor_0_resp_bits_tag),
		.io_requestor_0_resp_bits_data(dcacheArb_io_requestor_0_resp_bits_data),
		.io_requestor_0_resp_bits_replay(dcacheArb_io_requestor_0_resp_bits_replay),
		.io_requestor_0_resp_bits_has_data(dcacheArb_io_requestor_0_resp_bits_has_data),
		.io_requestor_0_resp_bits_data_word_bypass(dcacheArb_io_requestor_0_resp_bits_data_word_bypass),
		.io_requestor_0_replay_next(dcacheArb_io_requestor_0_replay_next),
		.io_requestor_0_s2_xcpt_ma_ld(dcacheArb_io_requestor_0_s2_xcpt_ma_ld),
		.io_requestor_0_s2_xcpt_ma_st(dcacheArb_io_requestor_0_s2_xcpt_ma_st),
		.io_requestor_0_s2_xcpt_pf_ld(dcacheArb_io_requestor_0_s2_xcpt_pf_ld),
		.io_requestor_0_s2_xcpt_pf_st(dcacheArb_io_requestor_0_s2_xcpt_pf_st),
		.io_requestor_0_s2_xcpt_ae_ld(dcacheArb_io_requestor_0_s2_xcpt_ae_ld),
		.io_requestor_0_s2_xcpt_ae_st(dcacheArb_io_requestor_0_s2_xcpt_ae_st),
		.io_requestor_0_ordered(dcacheArb_io_requestor_0_ordered),
		.io_requestor_0_perf_grant(dcacheArb_io_requestor_0_perf_grant),
		.io_requestor_1_req_ready(dcacheArb_io_requestor_1_req_ready),
		.io_requestor_1_req_valid(dcacheArb_io_requestor_1_req_valid),
		.io_requestor_1_req_bits_addr(dcacheArb_io_requestor_1_req_bits_addr),
		.io_requestor_1_req_bits_cmd(dcacheArb_io_requestor_1_req_bits_cmd),
		.io_requestor_1_req_bits_size(dcacheArb_io_requestor_1_req_bits_size),
		.io_requestor_1_s1_kill(dcacheArb_io_requestor_1_s1_kill),
		.io_requestor_1_s1_data_data(dcacheArb_io_requestor_1_s1_data_data),
		.io_requestor_1_s1_data_mask(dcacheArb_io_requestor_1_s1_data_mask),
		.io_requestor_1_s2_nack(dcacheArb_io_requestor_1_s2_nack),
		.io_requestor_1_resp_valid(dcacheArb_io_requestor_1_resp_valid),
		.io_requestor_1_resp_bits_data_raw(dcacheArb_io_requestor_1_resp_bits_data_raw),
		.io_mem_req_ready(dcacheArb_io_mem_req_ready),
		.io_mem_req_valid(dcacheArb_io_mem_req_valid),
		.io_mem_req_bits_addr(dcacheArb_io_mem_req_bits_addr),
		.io_mem_req_bits_tag(dcacheArb_io_mem_req_bits_tag),
		.io_mem_req_bits_cmd(dcacheArb_io_mem_req_bits_cmd),
		.io_mem_req_bits_size(dcacheArb_io_mem_req_bits_size),
		.io_mem_req_bits_signed(dcacheArb_io_mem_req_bits_signed),
		.io_mem_req_bits_dprv(dcacheArb_io_mem_req_bits_dprv),
		.io_mem_req_bits_no_xcpt(dcacheArb_io_mem_req_bits_no_xcpt),
		.io_mem_s1_kill(dcacheArb_io_mem_s1_kill),
		.io_mem_s1_data_data(dcacheArb_io_mem_s1_data_data),
		.io_mem_s1_data_mask(dcacheArb_io_mem_s1_data_mask),
		.io_mem_s2_nack(dcacheArb_io_mem_s2_nack),
		.io_mem_resp_valid(dcacheArb_io_mem_resp_valid),
		.io_mem_resp_bits_tag(dcacheArb_io_mem_resp_bits_tag),
		.io_mem_resp_bits_data(dcacheArb_io_mem_resp_bits_data),
		.io_mem_resp_bits_replay(dcacheArb_io_mem_resp_bits_replay),
		.io_mem_resp_bits_has_data(dcacheArb_io_mem_resp_bits_has_data),
		.io_mem_resp_bits_data_word_bypass(dcacheArb_io_mem_resp_bits_data_word_bypass),
		.io_mem_resp_bits_data_raw(dcacheArb_io_mem_resp_bits_data_raw),
		.io_mem_replay_next(dcacheArb_io_mem_replay_next),
		.io_mem_s2_xcpt_ma_ld(dcacheArb_io_mem_s2_xcpt_ma_ld),
		.io_mem_s2_xcpt_ma_st(dcacheArb_io_mem_s2_xcpt_ma_st),
		.io_mem_s2_xcpt_pf_ld(dcacheArb_io_mem_s2_xcpt_pf_ld),
		.io_mem_s2_xcpt_pf_st(dcacheArb_io_mem_s2_xcpt_pf_st),
		.io_mem_s2_xcpt_ae_ld(dcacheArb_io_mem_s2_xcpt_ae_ld),
		.io_mem_s2_xcpt_ae_st(dcacheArb_io_mem_s2_xcpt_ae_st),
		.io_mem_ordered(dcacheArb_io_mem_ordered),
		.io_mem_perf_grant(dcacheArb_io_mem_perf_grant)
	);
	PTW ptw(
		.clock(ptw_clock),
		.reset(ptw_reset),
		.io_requestor_0_status_debug(ptw_io_requestor_0_status_debug),
		.io_requestor_0_pmp_0_cfg_l(ptw_io_requestor_0_pmp_0_cfg_l),
		.io_requestor_0_pmp_0_cfg_a(ptw_io_requestor_0_pmp_0_cfg_a),
		.io_requestor_0_pmp_0_cfg_x(ptw_io_requestor_0_pmp_0_cfg_x),
		.io_requestor_0_pmp_0_cfg_w(ptw_io_requestor_0_pmp_0_cfg_w),
		.io_requestor_0_pmp_0_cfg_r(ptw_io_requestor_0_pmp_0_cfg_r),
		.io_requestor_0_pmp_0_addr(ptw_io_requestor_0_pmp_0_addr),
		.io_requestor_0_pmp_0_mask(ptw_io_requestor_0_pmp_0_mask),
		.io_requestor_0_pmp_1_cfg_l(ptw_io_requestor_0_pmp_1_cfg_l),
		.io_requestor_0_pmp_1_cfg_a(ptw_io_requestor_0_pmp_1_cfg_a),
		.io_requestor_0_pmp_1_cfg_x(ptw_io_requestor_0_pmp_1_cfg_x),
		.io_requestor_0_pmp_1_cfg_w(ptw_io_requestor_0_pmp_1_cfg_w),
		.io_requestor_0_pmp_1_cfg_r(ptw_io_requestor_0_pmp_1_cfg_r),
		.io_requestor_0_pmp_1_addr(ptw_io_requestor_0_pmp_1_addr),
		.io_requestor_0_pmp_1_mask(ptw_io_requestor_0_pmp_1_mask),
		.io_requestor_0_pmp_2_cfg_l(ptw_io_requestor_0_pmp_2_cfg_l),
		.io_requestor_0_pmp_2_cfg_a(ptw_io_requestor_0_pmp_2_cfg_a),
		.io_requestor_0_pmp_2_cfg_x(ptw_io_requestor_0_pmp_2_cfg_x),
		.io_requestor_0_pmp_2_cfg_w(ptw_io_requestor_0_pmp_2_cfg_w),
		.io_requestor_0_pmp_2_cfg_r(ptw_io_requestor_0_pmp_2_cfg_r),
		.io_requestor_0_pmp_2_addr(ptw_io_requestor_0_pmp_2_addr),
		.io_requestor_0_pmp_2_mask(ptw_io_requestor_0_pmp_2_mask),
		.io_requestor_0_pmp_3_cfg_l(ptw_io_requestor_0_pmp_3_cfg_l),
		.io_requestor_0_pmp_3_cfg_a(ptw_io_requestor_0_pmp_3_cfg_a),
		.io_requestor_0_pmp_3_cfg_x(ptw_io_requestor_0_pmp_3_cfg_x),
		.io_requestor_0_pmp_3_cfg_w(ptw_io_requestor_0_pmp_3_cfg_w),
		.io_requestor_0_pmp_3_cfg_r(ptw_io_requestor_0_pmp_3_cfg_r),
		.io_requestor_0_pmp_3_addr(ptw_io_requestor_0_pmp_3_addr),
		.io_requestor_0_pmp_3_mask(ptw_io_requestor_0_pmp_3_mask),
		.io_requestor_0_pmp_4_cfg_l(ptw_io_requestor_0_pmp_4_cfg_l),
		.io_requestor_0_pmp_4_cfg_a(ptw_io_requestor_0_pmp_4_cfg_a),
		.io_requestor_0_pmp_4_cfg_x(ptw_io_requestor_0_pmp_4_cfg_x),
		.io_requestor_0_pmp_4_cfg_w(ptw_io_requestor_0_pmp_4_cfg_w),
		.io_requestor_0_pmp_4_cfg_r(ptw_io_requestor_0_pmp_4_cfg_r),
		.io_requestor_0_pmp_4_addr(ptw_io_requestor_0_pmp_4_addr),
		.io_requestor_0_pmp_4_mask(ptw_io_requestor_0_pmp_4_mask),
		.io_requestor_0_pmp_5_cfg_l(ptw_io_requestor_0_pmp_5_cfg_l),
		.io_requestor_0_pmp_5_cfg_a(ptw_io_requestor_0_pmp_5_cfg_a),
		.io_requestor_0_pmp_5_cfg_x(ptw_io_requestor_0_pmp_5_cfg_x),
		.io_requestor_0_pmp_5_cfg_w(ptw_io_requestor_0_pmp_5_cfg_w),
		.io_requestor_0_pmp_5_cfg_r(ptw_io_requestor_0_pmp_5_cfg_r),
		.io_requestor_0_pmp_5_addr(ptw_io_requestor_0_pmp_5_addr),
		.io_requestor_0_pmp_5_mask(ptw_io_requestor_0_pmp_5_mask),
		.io_requestor_0_pmp_6_cfg_l(ptw_io_requestor_0_pmp_6_cfg_l),
		.io_requestor_0_pmp_6_cfg_a(ptw_io_requestor_0_pmp_6_cfg_a),
		.io_requestor_0_pmp_6_cfg_x(ptw_io_requestor_0_pmp_6_cfg_x),
		.io_requestor_0_pmp_6_cfg_w(ptw_io_requestor_0_pmp_6_cfg_w),
		.io_requestor_0_pmp_6_cfg_r(ptw_io_requestor_0_pmp_6_cfg_r),
		.io_requestor_0_pmp_6_addr(ptw_io_requestor_0_pmp_6_addr),
		.io_requestor_0_pmp_6_mask(ptw_io_requestor_0_pmp_6_mask),
		.io_requestor_0_pmp_7_cfg_l(ptw_io_requestor_0_pmp_7_cfg_l),
		.io_requestor_0_pmp_7_cfg_a(ptw_io_requestor_0_pmp_7_cfg_a),
		.io_requestor_0_pmp_7_cfg_x(ptw_io_requestor_0_pmp_7_cfg_x),
		.io_requestor_0_pmp_7_cfg_w(ptw_io_requestor_0_pmp_7_cfg_w),
		.io_requestor_0_pmp_7_cfg_r(ptw_io_requestor_0_pmp_7_cfg_r),
		.io_requestor_0_pmp_7_addr(ptw_io_requestor_0_pmp_7_addr),
		.io_requestor_0_pmp_7_mask(ptw_io_requestor_0_pmp_7_mask),
		.io_requestor_1_status_debug(ptw_io_requestor_1_status_debug),
		.io_requestor_1_pmp_0_cfg_l(ptw_io_requestor_1_pmp_0_cfg_l),
		.io_requestor_1_pmp_0_cfg_a(ptw_io_requestor_1_pmp_0_cfg_a),
		.io_requestor_1_pmp_0_cfg_x(ptw_io_requestor_1_pmp_0_cfg_x),
		.io_requestor_1_pmp_0_cfg_w(ptw_io_requestor_1_pmp_0_cfg_w),
		.io_requestor_1_pmp_0_cfg_r(ptw_io_requestor_1_pmp_0_cfg_r),
		.io_requestor_1_pmp_0_addr(ptw_io_requestor_1_pmp_0_addr),
		.io_requestor_1_pmp_0_mask(ptw_io_requestor_1_pmp_0_mask),
		.io_requestor_1_pmp_1_cfg_l(ptw_io_requestor_1_pmp_1_cfg_l),
		.io_requestor_1_pmp_1_cfg_a(ptw_io_requestor_1_pmp_1_cfg_a),
		.io_requestor_1_pmp_1_cfg_x(ptw_io_requestor_1_pmp_1_cfg_x),
		.io_requestor_1_pmp_1_cfg_w(ptw_io_requestor_1_pmp_1_cfg_w),
		.io_requestor_1_pmp_1_cfg_r(ptw_io_requestor_1_pmp_1_cfg_r),
		.io_requestor_1_pmp_1_addr(ptw_io_requestor_1_pmp_1_addr),
		.io_requestor_1_pmp_1_mask(ptw_io_requestor_1_pmp_1_mask),
		.io_requestor_1_pmp_2_cfg_l(ptw_io_requestor_1_pmp_2_cfg_l),
		.io_requestor_1_pmp_2_cfg_a(ptw_io_requestor_1_pmp_2_cfg_a),
		.io_requestor_1_pmp_2_cfg_x(ptw_io_requestor_1_pmp_2_cfg_x),
		.io_requestor_1_pmp_2_cfg_w(ptw_io_requestor_1_pmp_2_cfg_w),
		.io_requestor_1_pmp_2_cfg_r(ptw_io_requestor_1_pmp_2_cfg_r),
		.io_requestor_1_pmp_2_addr(ptw_io_requestor_1_pmp_2_addr),
		.io_requestor_1_pmp_2_mask(ptw_io_requestor_1_pmp_2_mask),
		.io_requestor_1_pmp_3_cfg_l(ptw_io_requestor_1_pmp_3_cfg_l),
		.io_requestor_1_pmp_3_cfg_a(ptw_io_requestor_1_pmp_3_cfg_a),
		.io_requestor_1_pmp_3_cfg_x(ptw_io_requestor_1_pmp_3_cfg_x),
		.io_requestor_1_pmp_3_cfg_w(ptw_io_requestor_1_pmp_3_cfg_w),
		.io_requestor_1_pmp_3_cfg_r(ptw_io_requestor_1_pmp_3_cfg_r),
		.io_requestor_1_pmp_3_addr(ptw_io_requestor_1_pmp_3_addr),
		.io_requestor_1_pmp_3_mask(ptw_io_requestor_1_pmp_3_mask),
		.io_requestor_1_pmp_4_cfg_l(ptw_io_requestor_1_pmp_4_cfg_l),
		.io_requestor_1_pmp_4_cfg_a(ptw_io_requestor_1_pmp_4_cfg_a),
		.io_requestor_1_pmp_4_cfg_x(ptw_io_requestor_1_pmp_4_cfg_x),
		.io_requestor_1_pmp_4_cfg_w(ptw_io_requestor_1_pmp_4_cfg_w),
		.io_requestor_1_pmp_4_cfg_r(ptw_io_requestor_1_pmp_4_cfg_r),
		.io_requestor_1_pmp_4_addr(ptw_io_requestor_1_pmp_4_addr),
		.io_requestor_1_pmp_4_mask(ptw_io_requestor_1_pmp_4_mask),
		.io_requestor_1_pmp_5_cfg_l(ptw_io_requestor_1_pmp_5_cfg_l),
		.io_requestor_1_pmp_5_cfg_a(ptw_io_requestor_1_pmp_5_cfg_a),
		.io_requestor_1_pmp_5_cfg_x(ptw_io_requestor_1_pmp_5_cfg_x),
		.io_requestor_1_pmp_5_cfg_w(ptw_io_requestor_1_pmp_5_cfg_w),
		.io_requestor_1_pmp_5_cfg_r(ptw_io_requestor_1_pmp_5_cfg_r),
		.io_requestor_1_pmp_5_addr(ptw_io_requestor_1_pmp_5_addr),
		.io_requestor_1_pmp_5_mask(ptw_io_requestor_1_pmp_5_mask),
		.io_requestor_1_pmp_6_cfg_l(ptw_io_requestor_1_pmp_6_cfg_l),
		.io_requestor_1_pmp_6_cfg_a(ptw_io_requestor_1_pmp_6_cfg_a),
		.io_requestor_1_pmp_6_cfg_x(ptw_io_requestor_1_pmp_6_cfg_x),
		.io_requestor_1_pmp_6_cfg_w(ptw_io_requestor_1_pmp_6_cfg_w),
		.io_requestor_1_pmp_6_cfg_r(ptw_io_requestor_1_pmp_6_cfg_r),
		.io_requestor_1_pmp_6_addr(ptw_io_requestor_1_pmp_6_addr),
		.io_requestor_1_pmp_6_mask(ptw_io_requestor_1_pmp_6_mask),
		.io_requestor_1_pmp_7_cfg_l(ptw_io_requestor_1_pmp_7_cfg_l),
		.io_requestor_1_pmp_7_cfg_a(ptw_io_requestor_1_pmp_7_cfg_a),
		.io_requestor_1_pmp_7_cfg_x(ptw_io_requestor_1_pmp_7_cfg_x),
		.io_requestor_1_pmp_7_cfg_w(ptw_io_requestor_1_pmp_7_cfg_w),
		.io_requestor_1_pmp_7_cfg_r(ptw_io_requestor_1_pmp_7_cfg_r),
		.io_requestor_1_pmp_7_addr(ptw_io_requestor_1_pmp_7_addr),
		.io_requestor_1_pmp_7_mask(ptw_io_requestor_1_pmp_7_mask),
		.io_requestor_1_customCSRs_csrs_0_value(ptw_io_requestor_1_customCSRs_csrs_0_value),
		.io_dpath_status_debug(ptw_io_dpath_status_debug),
		.io_dpath_pmp_0_cfg_l(ptw_io_dpath_pmp_0_cfg_l),
		.io_dpath_pmp_0_cfg_a(ptw_io_dpath_pmp_0_cfg_a),
		.io_dpath_pmp_0_cfg_x(ptw_io_dpath_pmp_0_cfg_x),
		.io_dpath_pmp_0_cfg_w(ptw_io_dpath_pmp_0_cfg_w),
		.io_dpath_pmp_0_cfg_r(ptw_io_dpath_pmp_0_cfg_r),
		.io_dpath_pmp_0_addr(ptw_io_dpath_pmp_0_addr),
		.io_dpath_pmp_0_mask(ptw_io_dpath_pmp_0_mask),
		.io_dpath_pmp_1_cfg_l(ptw_io_dpath_pmp_1_cfg_l),
		.io_dpath_pmp_1_cfg_a(ptw_io_dpath_pmp_1_cfg_a),
		.io_dpath_pmp_1_cfg_x(ptw_io_dpath_pmp_1_cfg_x),
		.io_dpath_pmp_1_cfg_w(ptw_io_dpath_pmp_1_cfg_w),
		.io_dpath_pmp_1_cfg_r(ptw_io_dpath_pmp_1_cfg_r),
		.io_dpath_pmp_1_addr(ptw_io_dpath_pmp_1_addr),
		.io_dpath_pmp_1_mask(ptw_io_dpath_pmp_1_mask),
		.io_dpath_pmp_2_cfg_l(ptw_io_dpath_pmp_2_cfg_l),
		.io_dpath_pmp_2_cfg_a(ptw_io_dpath_pmp_2_cfg_a),
		.io_dpath_pmp_2_cfg_x(ptw_io_dpath_pmp_2_cfg_x),
		.io_dpath_pmp_2_cfg_w(ptw_io_dpath_pmp_2_cfg_w),
		.io_dpath_pmp_2_cfg_r(ptw_io_dpath_pmp_2_cfg_r),
		.io_dpath_pmp_2_addr(ptw_io_dpath_pmp_2_addr),
		.io_dpath_pmp_2_mask(ptw_io_dpath_pmp_2_mask),
		.io_dpath_pmp_3_cfg_l(ptw_io_dpath_pmp_3_cfg_l),
		.io_dpath_pmp_3_cfg_a(ptw_io_dpath_pmp_3_cfg_a),
		.io_dpath_pmp_3_cfg_x(ptw_io_dpath_pmp_3_cfg_x),
		.io_dpath_pmp_3_cfg_w(ptw_io_dpath_pmp_3_cfg_w),
		.io_dpath_pmp_3_cfg_r(ptw_io_dpath_pmp_3_cfg_r),
		.io_dpath_pmp_3_addr(ptw_io_dpath_pmp_3_addr),
		.io_dpath_pmp_3_mask(ptw_io_dpath_pmp_3_mask),
		.io_dpath_pmp_4_cfg_l(ptw_io_dpath_pmp_4_cfg_l),
		.io_dpath_pmp_4_cfg_a(ptw_io_dpath_pmp_4_cfg_a),
		.io_dpath_pmp_4_cfg_x(ptw_io_dpath_pmp_4_cfg_x),
		.io_dpath_pmp_4_cfg_w(ptw_io_dpath_pmp_4_cfg_w),
		.io_dpath_pmp_4_cfg_r(ptw_io_dpath_pmp_4_cfg_r),
		.io_dpath_pmp_4_addr(ptw_io_dpath_pmp_4_addr),
		.io_dpath_pmp_4_mask(ptw_io_dpath_pmp_4_mask),
		.io_dpath_pmp_5_cfg_l(ptw_io_dpath_pmp_5_cfg_l),
		.io_dpath_pmp_5_cfg_a(ptw_io_dpath_pmp_5_cfg_a),
		.io_dpath_pmp_5_cfg_x(ptw_io_dpath_pmp_5_cfg_x),
		.io_dpath_pmp_5_cfg_w(ptw_io_dpath_pmp_5_cfg_w),
		.io_dpath_pmp_5_cfg_r(ptw_io_dpath_pmp_5_cfg_r),
		.io_dpath_pmp_5_addr(ptw_io_dpath_pmp_5_addr),
		.io_dpath_pmp_5_mask(ptw_io_dpath_pmp_5_mask),
		.io_dpath_pmp_6_cfg_l(ptw_io_dpath_pmp_6_cfg_l),
		.io_dpath_pmp_6_cfg_a(ptw_io_dpath_pmp_6_cfg_a),
		.io_dpath_pmp_6_cfg_x(ptw_io_dpath_pmp_6_cfg_x),
		.io_dpath_pmp_6_cfg_w(ptw_io_dpath_pmp_6_cfg_w),
		.io_dpath_pmp_6_cfg_r(ptw_io_dpath_pmp_6_cfg_r),
		.io_dpath_pmp_6_addr(ptw_io_dpath_pmp_6_addr),
		.io_dpath_pmp_6_mask(ptw_io_dpath_pmp_6_mask),
		.io_dpath_pmp_7_cfg_l(ptw_io_dpath_pmp_7_cfg_l),
		.io_dpath_pmp_7_cfg_a(ptw_io_dpath_pmp_7_cfg_a),
		.io_dpath_pmp_7_cfg_x(ptw_io_dpath_pmp_7_cfg_x),
		.io_dpath_pmp_7_cfg_w(ptw_io_dpath_pmp_7_cfg_w),
		.io_dpath_pmp_7_cfg_r(ptw_io_dpath_pmp_7_cfg_r),
		.io_dpath_pmp_7_addr(ptw_io_dpath_pmp_7_addr),
		.io_dpath_pmp_7_mask(ptw_io_dpath_pmp_7_mask),
		.io_dpath_perf_l2hit(ptw_io_dpath_perf_l2hit),
		.io_dpath_perf_pte_miss(ptw_io_dpath_perf_pte_miss),
		.io_dpath_perf_pte_hit(ptw_io_dpath_perf_pte_hit),
		.io_dpath_customCSRs_csrs_0_value(ptw_io_dpath_customCSRs_csrs_0_value)
	);
	Rocket core(
		.clock(core_clock),
		.reset(core_reset),
		.io_hartid(core_io_hartid),
		.io_interrupts_debug(core_io_interrupts_debug),
		.io_interrupts_mtip(core_io_interrupts_mtip),
		.io_interrupts_msip(core_io_interrupts_msip),
		.io_interrupts_meip(core_io_interrupts_meip),
		.io_imem_might_request(core_io_imem_might_request),
		.io_imem_req_valid(core_io_imem_req_valid),
		.io_imem_req_bits_pc(core_io_imem_req_bits_pc),
		.io_imem_req_bits_speculative(core_io_imem_req_bits_speculative),
		.io_imem_resp_ready(core_io_imem_resp_ready),
		.io_imem_resp_valid(core_io_imem_resp_valid),
		.io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
		.io_imem_resp_bits_data(core_io_imem_resp_bits_data),
		.io_imem_resp_bits_xcpt_ae_inst(core_io_imem_resp_bits_xcpt_ae_inst),
		.io_imem_resp_bits_replay(core_io_imem_resp_bits_replay),
		.io_imem_btb_update_valid(core_io_imem_btb_update_valid),
		.io_imem_bht_update_valid(core_io_imem_bht_update_valid),
		.io_imem_flush_icache(core_io_imem_flush_icache),
		.io_dmem_req_ready(core_io_dmem_req_ready),
		.io_dmem_req_valid(core_io_dmem_req_valid),
		.io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
		.io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
		.io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
		.io_dmem_req_bits_size(core_io_dmem_req_bits_size),
		.io_dmem_req_bits_signed(core_io_dmem_req_bits_signed),
		.io_dmem_req_bits_dv(core_io_dmem_req_bits_dv),
		.io_dmem_s1_kill(core_io_dmem_s1_kill),
		.io_dmem_s1_data_data(core_io_dmem_s1_data_data),
		.io_dmem_s2_nack(core_io_dmem_s2_nack),
		.io_dmem_resp_valid(core_io_dmem_resp_valid),
		.io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
		.io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
		.io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),
		.io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
		.io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),
		.io_dmem_replay_next(core_io_dmem_replay_next),
		.io_dmem_s2_xcpt_ma_ld(core_io_dmem_s2_xcpt_ma_ld),
		.io_dmem_s2_xcpt_ma_st(core_io_dmem_s2_xcpt_ma_st),
		.io_dmem_s2_xcpt_pf_ld(core_io_dmem_s2_xcpt_pf_ld),
		.io_dmem_s2_xcpt_pf_st(core_io_dmem_s2_xcpt_pf_st),
		.io_dmem_s2_xcpt_ae_ld(core_io_dmem_s2_xcpt_ae_ld),
		.io_dmem_s2_xcpt_ae_st(core_io_dmem_s2_xcpt_ae_st),
		.io_dmem_ordered(core_io_dmem_ordered),
		.io_dmem_perf_grant(core_io_dmem_perf_grant),
		.io_ptw_status_debug(core_io_ptw_status_debug),
		.io_ptw_pmp_0_cfg_l(core_io_ptw_pmp_0_cfg_l),
		.io_ptw_pmp_0_cfg_a(core_io_ptw_pmp_0_cfg_a),
		.io_ptw_pmp_0_cfg_x(core_io_ptw_pmp_0_cfg_x),
		.io_ptw_pmp_0_cfg_w(core_io_ptw_pmp_0_cfg_w),
		.io_ptw_pmp_0_cfg_r(core_io_ptw_pmp_0_cfg_r),
		.io_ptw_pmp_0_addr(core_io_ptw_pmp_0_addr),
		.io_ptw_pmp_0_mask(core_io_ptw_pmp_0_mask),
		.io_ptw_pmp_1_cfg_l(core_io_ptw_pmp_1_cfg_l),
		.io_ptw_pmp_1_cfg_a(core_io_ptw_pmp_1_cfg_a),
		.io_ptw_pmp_1_cfg_x(core_io_ptw_pmp_1_cfg_x),
		.io_ptw_pmp_1_cfg_w(core_io_ptw_pmp_1_cfg_w),
		.io_ptw_pmp_1_cfg_r(core_io_ptw_pmp_1_cfg_r),
		.io_ptw_pmp_1_addr(core_io_ptw_pmp_1_addr),
		.io_ptw_pmp_1_mask(core_io_ptw_pmp_1_mask),
		.io_ptw_pmp_2_cfg_l(core_io_ptw_pmp_2_cfg_l),
		.io_ptw_pmp_2_cfg_a(core_io_ptw_pmp_2_cfg_a),
		.io_ptw_pmp_2_cfg_x(core_io_ptw_pmp_2_cfg_x),
		.io_ptw_pmp_2_cfg_w(core_io_ptw_pmp_2_cfg_w),
		.io_ptw_pmp_2_cfg_r(core_io_ptw_pmp_2_cfg_r),
		.io_ptw_pmp_2_addr(core_io_ptw_pmp_2_addr),
		.io_ptw_pmp_2_mask(core_io_ptw_pmp_2_mask),
		.io_ptw_pmp_3_cfg_l(core_io_ptw_pmp_3_cfg_l),
		.io_ptw_pmp_3_cfg_a(core_io_ptw_pmp_3_cfg_a),
		.io_ptw_pmp_3_cfg_x(core_io_ptw_pmp_3_cfg_x),
		.io_ptw_pmp_3_cfg_w(core_io_ptw_pmp_3_cfg_w),
		.io_ptw_pmp_3_cfg_r(core_io_ptw_pmp_3_cfg_r),
		.io_ptw_pmp_3_addr(core_io_ptw_pmp_3_addr),
		.io_ptw_pmp_3_mask(core_io_ptw_pmp_3_mask),
		.io_ptw_pmp_4_cfg_l(core_io_ptw_pmp_4_cfg_l),
		.io_ptw_pmp_4_cfg_a(core_io_ptw_pmp_4_cfg_a),
		.io_ptw_pmp_4_cfg_x(core_io_ptw_pmp_4_cfg_x),
		.io_ptw_pmp_4_cfg_w(core_io_ptw_pmp_4_cfg_w),
		.io_ptw_pmp_4_cfg_r(core_io_ptw_pmp_4_cfg_r),
		.io_ptw_pmp_4_addr(core_io_ptw_pmp_4_addr),
		.io_ptw_pmp_4_mask(core_io_ptw_pmp_4_mask),
		.io_ptw_pmp_5_cfg_l(core_io_ptw_pmp_5_cfg_l),
		.io_ptw_pmp_5_cfg_a(core_io_ptw_pmp_5_cfg_a),
		.io_ptw_pmp_5_cfg_x(core_io_ptw_pmp_5_cfg_x),
		.io_ptw_pmp_5_cfg_w(core_io_ptw_pmp_5_cfg_w),
		.io_ptw_pmp_5_cfg_r(core_io_ptw_pmp_5_cfg_r),
		.io_ptw_pmp_5_addr(core_io_ptw_pmp_5_addr),
		.io_ptw_pmp_5_mask(core_io_ptw_pmp_5_mask),
		.io_ptw_pmp_6_cfg_l(core_io_ptw_pmp_6_cfg_l),
		.io_ptw_pmp_6_cfg_a(core_io_ptw_pmp_6_cfg_a),
		.io_ptw_pmp_6_cfg_x(core_io_ptw_pmp_6_cfg_x),
		.io_ptw_pmp_6_cfg_w(core_io_ptw_pmp_6_cfg_w),
		.io_ptw_pmp_6_cfg_r(core_io_ptw_pmp_6_cfg_r),
		.io_ptw_pmp_6_addr(core_io_ptw_pmp_6_addr),
		.io_ptw_pmp_6_mask(core_io_ptw_pmp_6_mask),
		.io_ptw_pmp_7_cfg_l(core_io_ptw_pmp_7_cfg_l),
		.io_ptw_pmp_7_cfg_a(core_io_ptw_pmp_7_cfg_a),
		.io_ptw_pmp_7_cfg_x(core_io_ptw_pmp_7_cfg_x),
		.io_ptw_pmp_7_cfg_w(core_io_ptw_pmp_7_cfg_w),
		.io_ptw_pmp_7_cfg_r(core_io_ptw_pmp_7_cfg_r),
		.io_ptw_pmp_7_addr(core_io_ptw_pmp_7_addr),
		.io_ptw_pmp_7_mask(core_io_ptw_pmp_7_mask),
		.io_ptw_customCSRs_csrs_0_value(core_io_ptw_customCSRs_csrs_0_value),
		.io_wfi(core_io_wfi)
	);
	assign auto_slave_in_a_ready = tlSlaveXbar_auto_in_a_ready;
	assign auto_slave_in_d_valid = tlSlaveXbar_auto_in_d_valid;
	assign auto_slave_in_d_bits_opcode = tlSlaveXbar_auto_in_d_bits_opcode;
	assign auto_slave_in_d_bits_size = tlSlaveXbar_auto_in_d_bits_size;
	assign auto_slave_in_d_bits_source = tlSlaveXbar_auto_in_d_bits_source;
	assign auto_slave_in_d_bits_data = tlSlaveXbar_auto_in_d_bits_data;
	assign auto_wfi_out_0 = bundleOut_0_0_REG;
	assign auto_tl_other_masters_out_a_valid = tlMasterXbar_auto_out_a_valid;
	assign auto_tl_other_masters_out_a_bits_opcode = tlMasterXbar_auto_out_a_bits_opcode;
	assign auto_tl_other_masters_out_a_bits_param = tlMasterXbar_auto_out_a_bits_param;
	assign auto_tl_other_masters_out_a_bits_size = tlMasterXbar_auto_out_a_bits_size;
	assign auto_tl_other_masters_out_a_bits_source = tlMasterXbar_auto_out_a_bits_source;
	assign auto_tl_other_masters_out_a_bits_address = tlMasterXbar_auto_out_a_bits_address;
	assign auto_tl_other_masters_out_a_bits_mask = tlMasterXbar_auto_out_a_bits_mask;
	assign auto_tl_other_masters_out_a_bits_data = tlMasterXbar_auto_out_a_bits_data;
	assign auto_tl_other_masters_out_d_ready = tlMasterXbar_auto_out_d_ready;
	assign tlMasterXbar_clock = clock;
	assign tlMasterXbar_reset = reset;
	assign tlMasterXbar_auto_in_1_a_valid = frontend_auto_icache_master_out_a_valid;
	assign tlMasterXbar_auto_in_1_a_bits_address = frontend_auto_icache_master_out_a_bits_address;
	assign tlMasterXbar_auto_in_0_a_valid = dcache_auto_out_a_valid;
	assign tlMasterXbar_auto_in_0_a_bits_opcode = dcache_auto_out_a_bits_opcode;
	assign tlMasterXbar_auto_in_0_a_bits_param = dcache_auto_out_a_bits_param;
	assign tlMasterXbar_auto_in_0_a_bits_size = dcache_auto_out_a_bits_size;
	assign tlMasterXbar_auto_in_0_a_bits_address = dcache_auto_out_a_bits_address;
	assign tlMasterXbar_auto_in_0_a_bits_mask = dcache_auto_out_a_bits_mask;
	assign tlMasterXbar_auto_in_0_a_bits_data = dcache_auto_out_a_bits_data;
	assign tlMasterXbar_auto_in_0_d_ready = dcache_auto_out_d_ready;
	assign tlMasterXbar_auto_out_a_ready = auto_tl_other_masters_out_a_ready;
	assign tlMasterXbar_auto_out_d_valid = auto_tl_other_masters_out_d_valid;
	assign tlMasterXbar_auto_out_d_bits_opcode = auto_tl_other_masters_out_d_bits_opcode;
	assign tlMasterXbar_auto_out_d_bits_param = auto_tl_other_masters_out_d_bits_param;
	assign tlMasterXbar_auto_out_d_bits_size = auto_tl_other_masters_out_d_bits_size;
	assign tlMasterXbar_auto_out_d_bits_source = auto_tl_other_masters_out_d_bits_source;
	assign tlMasterXbar_auto_out_d_bits_sink = auto_tl_other_masters_out_d_bits_sink;
	assign tlMasterXbar_auto_out_d_bits_denied = auto_tl_other_masters_out_d_bits_denied;
	assign tlMasterXbar_auto_out_d_bits_data = auto_tl_other_masters_out_d_bits_data;
	assign tlMasterXbar_auto_out_d_bits_corrupt = auto_tl_other_masters_out_d_bits_corrupt;
	assign tlSlaveXbar_auto_in_a_valid = auto_slave_in_a_valid;
	assign tlSlaveXbar_auto_in_a_bits_opcode = auto_slave_in_a_bits_opcode;
	assign tlSlaveXbar_auto_in_a_bits_param = auto_slave_in_a_bits_param;
	assign tlSlaveXbar_auto_in_a_bits_size = auto_slave_in_a_bits_size;
	assign tlSlaveXbar_auto_in_a_bits_source = auto_slave_in_a_bits_source;
	assign tlSlaveXbar_auto_in_a_bits_address = auto_slave_in_a_bits_address;
	assign tlSlaveXbar_auto_in_a_bits_mask = auto_slave_in_a_bits_mask;
	assign tlSlaveXbar_auto_in_a_bits_data = auto_slave_in_a_bits_data;
	assign tlSlaveXbar_auto_in_d_ready = auto_slave_in_d_ready;
	assign tlSlaveXbar_auto_out_a_ready = fragmenter_1_auto_in_a_ready;
	assign tlSlaveXbar_auto_out_d_valid = fragmenter_1_auto_in_d_valid;
	assign tlSlaveXbar_auto_out_d_bits_opcode = fragmenter_1_auto_in_d_bits_opcode;
	assign tlSlaveXbar_auto_out_d_bits_size = fragmenter_1_auto_in_d_bits_size;
	assign tlSlaveXbar_auto_out_d_bits_source = fragmenter_1_auto_in_d_bits_source;
	assign tlSlaveXbar_auto_out_d_bits_data = fragmenter_1_auto_in_d_bits_data;
	assign intXbar_auto_int_in_2_0 = auto_int_local_in_2_0;
	assign intXbar_auto_int_in_1_0 = auto_int_local_in_1_0;
	assign intXbar_auto_int_in_1_1 = auto_int_local_in_1_1;
	assign intXbar_auto_int_in_0_0 = auto_int_local_in_0_0;
	assign broadcast_auto_in = auto_hartid_in;
	assign dcache_clock = clock;
	assign dcache_reset = reset;
	assign dcache_auto_out_a_ready = tlMasterXbar_auto_in_0_a_ready;
	assign dcache_auto_out_d_valid = tlMasterXbar_auto_in_0_d_valid;
	assign dcache_auto_out_d_bits_opcode = tlMasterXbar_auto_in_0_d_bits_opcode;
	assign dcache_auto_out_d_bits_size = tlMasterXbar_auto_in_0_d_bits_size;
	assign dcache_auto_out_d_bits_denied = tlMasterXbar_auto_in_0_d_bits_denied;
	assign dcache_auto_out_d_bits_data = tlMasterXbar_auto_in_0_d_bits_data;
	assign dcache_io_cpu_req_valid = dcacheArb_io_mem_req_valid;
	assign dcache_io_cpu_req_bits_addr = dcacheArb_io_mem_req_bits_addr;
	assign dcache_io_cpu_req_bits_tag = dcacheArb_io_mem_req_bits_tag;
	assign dcache_io_cpu_req_bits_cmd = dcacheArb_io_mem_req_bits_cmd;
	assign dcache_io_cpu_req_bits_size = dcacheArb_io_mem_req_bits_size;
	assign dcache_io_cpu_req_bits_signed = dcacheArb_io_mem_req_bits_signed;
	assign dcache_io_cpu_req_bits_dprv = dcacheArb_io_mem_req_bits_dprv;
	assign dcache_io_cpu_req_bits_no_xcpt = dcacheArb_io_mem_req_bits_no_xcpt;
	assign dcache_io_cpu_s1_kill = dcacheArb_io_mem_s1_kill;
	assign dcache_io_cpu_s1_data_data = dcacheArb_io_mem_s1_data_data;
	assign dcache_io_cpu_s1_data_mask = dcacheArb_io_mem_s1_data_mask;
	assign dcache_io_ptw_status_debug = ptw_io_requestor_0_status_debug;
	assign dcache_io_ptw_pmp_0_cfg_l = ptw_io_requestor_0_pmp_0_cfg_l;
	assign dcache_io_ptw_pmp_0_cfg_a = ptw_io_requestor_0_pmp_0_cfg_a;
	assign dcache_io_ptw_pmp_0_cfg_x = ptw_io_requestor_0_pmp_0_cfg_x;
	assign dcache_io_ptw_pmp_0_cfg_w = ptw_io_requestor_0_pmp_0_cfg_w;
	assign dcache_io_ptw_pmp_0_cfg_r = ptw_io_requestor_0_pmp_0_cfg_r;
	assign dcache_io_ptw_pmp_0_addr = ptw_io_requestor_0_pmp_0_addr;
	assign dcache_io_ptw_pmp_0_mask = ptw_io_requestor_0_pmp_0_mask;
	assign dcache_io_ptw_pmp_1_cfg_l = ptw_io_requestor_0_pmp_1_cfg_l;
	assign dcache_io_ptw_pmp_1_cfg_a = ptw_io_requestor_0_pmp_1_cfg_a;
	assign dcache_io_ptw_pmp_1_cfg_x = ptw_io_requestor_0_pmp_1_cfg_x;
	assign dcache_io_ptw_pmp_1_cfg_w = ptw_io_requestor_0_pmp_1_cfg_w;
	assign dcache_io_ptw_pmp_1_cfg_r = ptw_io_requestor_0_pmp_1_cfg_r;
	assign dcache_io_ptw_pmp_1_addr = ptw_io_requestor_0_pmp_1_addr;
	assign dcache_io_ptw_pmp_1_mask = ptw_io_requestor_0_pmp_1_mask;
	assign dcache_io_ptw_pmp_2_cfg_l = ptw_io_requestor_0_pmp_2_cfg_l;
	assign dcache_io_ptw_pmp_2_cfg_a = ptw_io_requestor_0_pmp_2_cfg_a;
	assign dcache_io_ptw_pmp_2_cfg_x = ptw_io_requestor_0_pmp_2_cfg_x;
	assign dcache_io_ptw_pmp_2_cfg_w = ptw_io_requestor_0_pmp_2_cfg_w;
	assign dcache_io_ptw_pmp_2_cfg_r = ptw_io_requestor_0_pmp_2_cfg_r;
	assign dcache_io_ptw_pmp_2_addr = ptw_io_requestor_0_pmp_2_addr;
	assign dcache_io_ptw_pmp_2_mask = ptw_io_requestor_0_pmp_2_mask;
	assign dcache_io_ptw_pmp_3_cfg_l = ptw_io_requestor_0_pmp_3_cfg_l;
	assign dcache_io_ptw_pmp_3_cfg_a = ptw_io_requestor_0_pmp_3_cfg_a;
	assign dcache_io_ptw_pmp_3_cfg_x = ptw_io_requestor_0_pmp_3_cfg_x;
	assign dcache_io_ptw_pmp_3_cfg_w = ptw_io_requestor_0_pmp_3_cfg_w;
	assign dcache_io_ptw_pmp_3_cfg_r = ptw_io_requestor_0_pmp_3_cfg_r;
	assign dcache_io_ptw_pmp_3_addr = ptw_io_requestor_0_pmp_3_addr;
	assign dcache_io_ptw_pmp_3_mask = ptw_io_requestor_0_pmp_3_mask;
	assign dcache_io_ptw_pmp_4_cfg_l = ptw_io_requestor_0_pmp_4_cfg_l;
	assign dcache_io_ptw_pmp_4_cfg_a = ptw_io_requestor_0_pmp_4_cfg_a;
	assign dcache_io_ptw_pmp_4_cfg_x = ptw_io_requestor_0_pmp_4_cfg_x;
	assign dcache_io_ptw_pmp_4_cfg_w = ptw_io_requestor_0_pmp_4_cfg_w;
	assign dcache_io_ptw_pmp_4_cfg_r = ptw_io_requestor_0_pmp_4_cfg_r;
	assign dcache_io_ptw_pmp_4_addr = ptw_io_requestor_0_pmp_4_addr;
	assign dcache_io_ptw_pmp_4_mask = ptw_io_requestor_0_pmp_4_mask;
	assign dcache_io_ptw_pmp_5_cfg_l = ptw_io_requestor_0_pmp_5_cfg_l;
	assign dcache_io_ptw_pmp_5_cfg_a = ptw_io_requestor_0_pmp_5_cfg_a;
	assign dcache_io_ptw_pmp_5_cfg_x = ptw_io_requestor_0_pmp_5_cfg_x;
	assign dcache_io_ptw_pmp_5_cfg_w = ptw_io_requestor_0_pmp_5_cfg_w;
	assign dcache_io_ptw_pmp_5_cfg_r = ptw_io_requestor_0_pmp_5_cfg_r;
	assign dcache_io_ptw_pmp_5_addr = ptw_io_requestor_0_pmp_5_addr;
	assign dcache_io_ptw_pmp_5_mask = ptw_io_requestor_0_pmp_5_mask;
	assign dcache_io_ptw_pmp_6_cfg_l = ptw_io_requestor_0_pmp_6_cfg_l;
	assign dcache_io_ptw_pmp_6_cfg_a = ptw_io_requestor_0_pmp_6_cfg_a;
	assign dcache_io_ptw_pmp_6_cfg_x = ptw_io_requestor_0_pmp_6_cfg_x;
	assign dcache_io_ptw_pmp_6_cfg_w = ptw_io_requestor_0_pmp_6_cfg_w;
	assign dcache_io_ptw_pmp_6_cfg_r = ptw_io_requestor_0_pmp_6_cfg_r;
	assign dcache_io_ptw_pmp_6_addr = ptw_io_requestor_0_pmp_6_addr;
	assign dcache_io_ptw_pmp_6_mask = ptw_io_requestor_0_pmp_6_mask;
	assign dcache_io_ptw_pmp_7_cfg_l = ptw_io_requestor_0_pmp_7_cfg_l;
	assign dcache_io_ptw_pmp_7_cfg_a = ptw_io_requestor_0_pmp_7_cfg_a;
	assign dcache_io_ptw_pmp_7_cfg_x = ptw_io_requestor_0_pmp_7_cfg_x;
	assign dcache_io_ptw_pmp_7_cfg_w = ptw_io_requestor_0_pmp_7_cfg_w;
	assign dcache_io_ptw_pmp_7_cfg_r = ptw_io_requestor_0_pmp_7_cfg_r;
	assign dcache_io_ptw_pmp_7_addr = ptw_io_requestor_0_pmp_7_addr;
	assign dcache_io_ptw_pmp_7_mask = ptw_io_requestor_0_pmp_7_mask;
	assign frontend_clock = clock;
	assign frontend_reset = reset;
	assign frontend_auto_icache_master_out_a_ready = tlMasterXbar_auto_in_1_a_ready;
	assign frontend_auto_icache_master_out_d_valid = tlMasterXbar_auto_in_1_d_valid;
	assign frontend_auto_icache_master_out_d_bits_opcode = tlMasterXbar_auto_in_1_d_bits_opcode;
	assign frontend_auto_icache_master_out_d_bits_size = tlMasterXbar_auto_in_1_d_bits_size;
	assign frontend_auto_icache_master_out_d_bits_data = tlMasterXbar_auto_in_1_d_bits_data;
	assign frontend_auto_icache_master_out_d_bits_corrupt = tlMasterXbar_auto_in_1_d_bits_corrupt;
	assign frontend_io_cpu_might_request = core_io_imem_might_request;
	assign frontend_io_cpu_req_valid = core_io_imem_req_valid;
	assign frontend_io_cpu_req_bits_pc = core_io_imem_req_bits_pc;
	assign frontend_io_cpu_req_bits_speculative = core_io_imem_req_bits_speculative;
	assign frontend_io_cpu_resp_ready = core_io_imem_resp_ready;
	assign frontend_io_cpu_btb_update_valid = core_io_imem_btb_update_valid;
	assign frontend_io_cpu_bht_update_valid = core_io_imem_bht_update_valid;
	assign frontend_io_cpu_flush_icache = core_io_imem_flush_icache;
	assign frontend_io_ptw_status_debug = ptw_io_requestor_1_status_debug;
	assign frontend_io_ptw_pmp_0_cfg_l = ptw_io_requestor_1_pmp_0_cfg_l;
	assign frontend_io_ptw_pmp_0_cfg_a = ptw_io_requestor_1_pmp_0_cfg_a;
	assign frontend_io_ptw_pmp_0_cfg_x = ptw_io_requestor_1_pmp_0_cfg_x;
	assign frontend_io_ptw_pmp_0_cfg_w = ptw_io_requestor_1_pmp_0_cfg_w;
	assign frontend_io_ptw_pmp_0_cfg_r = ptw_io_requestor_1_pmp_0_cfg_r;
	assign frontend_io_ptw_pmp_0_addr = ptw_io_requestor_1_pmp_0_addr;
	assign frontend_io_ptw_pmp_0_mask = ptw_io_requestor_1_pmp_0_mask;
	assign frontend_io_ptw_pmp_1_cfg_l = ptw_io_requestor_1_pmp_1_cfg_l;
	assign frontend_io_ptw_pmp_1_cfg_a = ptw_io_requestor_1_pmp_1_cfg_a;
	assign frontend_io_ptw_pmp_1_cfg_x = ptw_io_requestor_1_pmp_1_cfg_x;
	assign frontend_io_ptw_pmp_1_cfg_w = ptw_io_requestor_1_pmp_1_cfg_w;
	assign frontend_io_ptw_pmp_1_cfg_r = ptw_io_requestor_1_pmp_1_cfg_r;
	assign frontend_io_ptw_pmp_1_addr = ptw_io_requestor_1_pmp_1_addr;
	assign frontend_io_ptw_pmp_1_mask = ptw_io_requestor_1_pmp_1_mask;
	assign frontend_io_ptw_pmp_2_cfg_l = ptw_io_requestor_1_pmp_2_cfg_l;
	assign frontend_io_ptw_pmp_2_cfg_a = ptw_io_requestor_1_pmp_2_cfg_a;
	assign frontend_io_ptw_pmp_2_cfg_x = ptw_io_requestor_1_pmp_2_cfg_x;
	assign frontend_io_ptw_pmp_2_cfg_w = ptw_io_requestor_1_pmp_2_cfg_w;
	assign frontend_io_ptw_pmp_2_cfg_r = ptw_io_requestor_1_pmp_2_cfg_r;
	assign frontend_io_ptw_pmp_2_addr = ptw_io_requestor_1_pmp_2_addr;
	assign frontend_io_ptw_pmp_2_mask = ptw_io_requestor_1_pmp_2_mask;
	assign frontend_io_ptw_pmp_3_cfg_l = ptw_io_requestor_1_pmp_3_cfg_l;
	assign frontend_io_ptw_pmp_3_cfg_a = ptw_io_requestor_1_pmp_3_cfg_a;
	assign frontend_io_ptw_pmp_3_cfg_x = ptw_io_requestor_1_pmp_3_cfg_x;
	assign frontend_io_ptw_pmp_3_cfg_w = ptw_io_requestor_1_pmp_3_cfg_w;
	assign frontend_io_ptw_pmp_3_cfg_r = ptw_io_requestor_1_pmp_3_cfg_r;
	assign frontend_io_ptw_pmp_3_addr = ptw_io_requestor_1_pmp_3_addr;
	assign frontend_io_ptw_pmp_3_mask = ptw_io_requestor_1_pmp_3_mask;
	assign frontend_io_ptw_pmp_4_cfg_l = ptw_io_requestor_1_pmp_4_cfg_l;
	assign frontend_io_ptw_pmp_4_cfg_a = ptw_io_requestor_1_pmp_4_cfg_a;
	assign frontend_io_ptw_pmp_4_cfg_x = ptw_io_requestor_1_pmp_4_cfg_x;
	assign frontend_io_ptw_pmp_4_cfg_w = ptw_io_requestor_1_pmp_4_cfg_w;
	assign frontend_io_ptw_pmp_4_cfg_r = ptw_io_requestor_1_pmp_4_cfg_r;
	assign frontend_io_ptw_pmp_4_addr = ptw_io_requestor_1_pmp_4_addr;
	assign frontend_io_ptw_pmp_4_mask = ptw_io_requestor_1_pmp_4_mask;
	assign frontend_io_ptw_pmp_5_cfg_l = ptw_io_requestor_1_pmp_5_cfg_l;
	assign frontend_io_ptw_pmp_5_cfg_a = ptw_io_requestor_1_pmp_5_cfg_a;
	assign frontend_io_ptw_pmp_5_cfg_x = ptw_io_requestor_1_pmp_5_cfg_x;
	assign frontend_io_ptw_pmp_5_cfg_w = ptw_io_requestor_1_pmp_5_cfg_w;
	assign frontend_io_ptw_pmp_5_cfg_r = ptw_io_requestor_1_pmp_5_cfg_r;
	assign frontend_io_ptw_pmp_5_addr = ptw_io_requestor_1_pmp_5_addr;
	assign frontend_io_ptw_pmp_5_mask = ptw_io_requestor_1_pmp_5_mask;
	assign frontend_io_ptw_pmp_6_cfg_l = ptw_io_requestor_1_pmp_6_cfg_l;
	assign frontend_io_ptw_pmp_6_cfg_a = ptw_io_requestor_1_pmp_6_cfg_a;
	assign frontend_io_ptw_pmp_6_cfg_x = ptw_io_requestor_1_pmp_6_cfg_x;
	assign frontend_io_ptw_pmp_6_cfg_w = ptw_io_requestor_1_pmp_6_cfg_w;
	assign frontend_io_ptw_pmp_6_cfg_r = ptw_io_requestor_1_pmp_6_cfg_r;
	assign frontend_io_ptw_pmp_6_addr = ptw_io_requestor_1_pmp_6_addr;
	assign frontend_io_ptw_pmp_6_mask = ptw_io_requestor_1_pmp_6_mask;
	assign frontend_io_ptw_pmp_7_cfg_l = ptw_io_requestor_1_pmp_7_cfg_l;
	assign frontend_io_ptw_pmp_7_cfg_a = ptw_io_requestor_1_pmp_7_cfg_a;
	assign frontend_io_ptw_pmp_7_cfg_x = ptw_io_requestor_1_pmp_7_cfg_x;
	assign frontend_io_ptw_pmp_7_cfg_w = ptw_io_requestor_1_pmp_7_cfg_w;
	assign frontend_io_ptw_pmp_7_cfg_r = ptw_io_requestor_1_pmp_7_cfg_r;
	assign frontend_io_ptw_pmp_7_addr = ptw_io_requestor_1_pmp_7_addr;
	assign frontend_io_ptw_pmp_7_mask = ptw_io_requestor_1_pmp_7_mask;
	assign frontend_io_ptw_customCSRs_csrs_0_value = ptw_io_requestor_1_customCSRs_csrs_0_value;
	assign dtim_adapter_clock = clock;
	assign dtim_adapter_reset = reset;
	assign dtim_adapter_auto_in_a_valid = fragmenter_1_auto_out_a_valid;
	assign dtim_adapter_auto_in_a_bits_opcode = fragmenter_1_auto_out_a_bits_opcode;
	assign dtim_adapter_auto_in_a_bits_param = fragmenter_1_auto_out_a_bits_param;
	assign dtim_adapter_auto_in_a_bits_size = fragmenter_1_auto_out_a_bits_size;
	assign dtim_adapter_auto_in_a_bits_source = fragmenter_1_auto_out_a_bits_source;
	assign dtim_adapter_auto_in_a_bits_address = fragmenter_1_auto_out_a_bits_address;
	assign dtim_adapter_auto_in_a_bits_mask = fragmenter_1_auto_out_a_bits_mask;
	assign dtim_adapter_auto_in_a_bits_data = fragmenter_1_auto_out_a_bits_data;
	assign dtim_adapter_auto_in_d_ready = fragmenter_1_auto_out_d_ready;
	assign dtim_adapter_io_dmem_req_ready = dcacheArb_io_requestor_1_req_ready;
	assign dtim_adapter_io_dmem_s2_nack = dcacheArb_io_requestor_1_s2_nack;
	assign dtim_adapter_io_dmem_resp_valid = dcacheArb_io_requestor_1_resp_valid;
	assign dtim_adapter_io_dmem_resp_bits_data_raw = dcacheArb_io_requestor_1_resp_bits_data_raw;
	assign fragmenter_1_clock = clock;
	assign fragmenter_1_reset = reset;
	assign fragmenter_1_auto_in_a_valid = tlSlaveXbar_auto_out_a_valid;
	assign fragmenter_1_auto_in_a_bits_opcode = tlSlaveXbar_auto_out_a_bits_opcode;
	assign fragmenter_1_auto_in_a_bits_param = tlSlaveXbar_auto_out_a_bits_param;
	assign fragmenter_1_auto_in_a_bits_size = tlSlaveXbar_auto_out_a_bits_size;
	assign fragmenter_1_auto_in_a_bits_source = tlSlaveXbar_auto_out_a_bits_source;
	assign fragmenter_1_auto_in_a_bits_address = tlSlaveXbar_auto_out_a_bits_address;
	assign fragmenter_1_auto_in_a_bits_mask = tlSlaveXbar_auto_out_a_bits_mask;
	assign fragmenter_1_auto_in_a_bits_data = tlSlaveXbar_auto_out_a_bits_data;
	assign fragmenter_1_auto_in_d_ready = tlSlaveXbar_auto_out_d_ready;
	assign fragmenter_1_auto_out_a_ready = dtim_adapter_auto_in_a_ready;
	assign fragmenter_1_auto_out_d_valid = dtim_adapter_auto_in_d_valid;
	assign fragmenter_1_auto_out_d_bits_opcode = dtim_adapter_auto_in_d_bits_opcode;
	assign fragmenter_1_auto_out_d_bits_size = dtim_adapter_auto_in_d_bits_size;
	assign fragmenter_1_auto_out_d_bits_source = dtim_adapter_auto_in_d_bits_source;
	assign fragmenter_1_auto_out_d_bits_data = dtim_adapter_auto_in_d_bits_data;
	assign dcacheArb_clock = clock;
	assign dcacheArb_io_requestor_0_req_valid = core_io_dmem_req_valid;
	assign dcacheArb_io_requestor_0_req_bits_addr = core_io_dmem_req_bits_addr;
	assign dcacheArb_io_requestor_0_req_bits_tag = core_io_dmem_req_bits_tag;
	assign dcacheArb_io_requestor_0_req_bits_cmd = core_io_dmem_req_bits_cmd;
	assign dcacheArb_io_requestor_0_req_bits_size = core_io_dmem_req_bits_size;
	assign dcacheArb_io_requestor_0_req_bits_signed = core_io_dmem_req_bits_signed;
	assign dcacheArb_io_requestor_0_s1_kill = core_io_dmem_s1_kill;
	assign dcacheArb_io_requestor_0_s1_data_data = core_io_dmem_s1_data_data;
	assign dcacheArb_io_requestor_1_req_valid = dtim_adapter_io_dmem_req_valid;
	assign dcacheArb_io_requestor_1_req_bits_addr = dtim_adapter_io_dmem_req_bits_addr;
	assign dcacheArb_io_requestor_1_req_bits_cmd = dtim_adapter_io_dmem_req_bits_cmd;
	assign dcacheArb_io_requestor_1_req_bits_size = dtim_adapter_io_dmem_req_bits_size;
	assign dcacheArb_io_requestor_1_s1_kill = dtim_adapter_io_dmem_s1_kill;
	assign dcacheArb_io_requestor_1_s1_data_data = dtim_adapter_io_dmem_s1_data_data;
	assign dcacheArb_io_requestor_1_s1_data_mask = dtim_adapter_io_dmem_s1_data_mask;
	assign dcacheArb_io_mem_req_ready = dcache_io_cpu_req_ready;
	assign dcacheArb_io_mem_s2_nack = dcache_io_cpu_s2_nack;
	assign dcacheArb_io_mem_resp_valid = dcache_io_cpu_resp_valid;
	assign dcacheArb_io_mem_resp_bits_tag = dcache_io_cpu_resp_bits_tag;
	assign dcacheArb_io_mem_resp_bits_data = dcache_io_cpu_resp_bits_data;
	assign dcacheArb_io_mem_resp_bits_replay = dcache_io_cpu_resp_bits_replay;
	assign dcacheArb_io_mem_resp_bits_has_data = dcache_io_cpu_resp_bits_has_data;
	assign dcacheArb_io_mem_resp_bits_data_word_bypass = dcache_io_cpu_resp_bits_data_word_bypass;
	assign dcacheArb_io_mem_resp_bits_data_raw = dcache_io_cpu_resp_bits_data_raw;
	assign dcacheArb_io_mem_replay_next = dcache_io_cpu_replay_next;
	assign dcacheArb_io_mem_s2_xcpt_ma_ld = dcache_io_cpu_s2_xcpt_ma_ld;
	assign dcacheArb_io_mem_s2_xcpt_ma_st = dcache_io_cpu_s2_xcpt_ma_st;
	assign dcacheArb_io_mem_s2_xcpt_pf_ld = dcache_io_cpu_s2_xcpt_pf_ld;
	assign dcacheArb_io_mem_s2_xcpt_pf_st = dcache_io_cpu_s2_xcpt_pf_st;
	assign dcacheArb_io_mem_s2_xcpt_ae_ld = dcache_io_cpu_s2_xcpt_ae_ld;
	assign dcacheArb_io_mem_s2_xcpt_ae_st = dcache_io_cpu_s2_xcpt_ae_st;
	assign dcacheArb_io_mem_ordered = dcache_io_cpu_ordered;
	assign dcacheArb_io_mem_perf_grant = dcache_io_cpu_perf_grant;
	assign ptw_clock = clock;
	assign ptw_reset = reset;
	assign ptw_io_dpath_status_debug = core_io_ptw_status_debug;
	assign ptw_io_dpath_pmp_0_cfg_l = core_io_ptw_pmp_0_cfg_l;
	assign ptw_io_dpath_pmp_0_cfg_a = core_io_ptw_pmp_0_cfg_a;
	assign ptw_io_dpath_pmp_0_cfg_x = core_io_ptw_pmp_0_cfg_x;
	assign ptw_io_dpath_pmp_0_cfg_w = core_io_ptw_pmp_0_cfg_w;
	assign ptw_io_dpath_pmp_0_cfg_r = core_io_ptw_pmp_0_cfg_r;
	assign ptw_io_dpath_pmp_0_addr = core_io_ptw_pmp_0_addr;
	assign ptw_io_dpath_pmp_0_mask = core_io_ptw_pmp_0_mask;
	assign ptw_io_dpath_pmp_1_cfg_l = core_io_ptw_pmp_1_cfg_l;
	assign ptw_io_dpath_pmp_1_cfg_a = core_io_ptw_pmp_1_cfg_a;
	assign ptw_io_dpath_pmp_1_cfg_x = core_io_ptw_pmp_1_cfg_x;
	assign ptw_io_dpath_pmp_1_cfg_w = core_io_ptw_pmp_1_cfg_w;
	assign ptw_io_dpath_pmp_1_cfg_r = core_io_ptw_pmp_1_cfg_r;
	assign ptw_io_dpath_pmp_1_addr = core_io_ptw_pmp_1_addr;
	assign ptw_io_dpath_pmp_1_mask = core_io_ptw_pmp_1_mask;
	assign ptw_io_dpath_pmp_2_cfg_l = core_io_ptw_pmp_2_cfg_l;
	assign ptw_io_dpath_pmp_2_cfg_a = core_io_ptw_pmp_2_cfg_a;
	assign ptw_io_dpath_pmp_2_cfg_x = core_io_ptw_pmp_2_cfg_x;
	assign ptw_io_dpath_pmp_2_cfg_w = core_io_ptw_pmp_2_cfg_w;
	assign ptw_io_dpath_pmp_2_cfg_r = core_io_ptw_pmp_2_cfg_r;
	assign ptw_io_dpath_pmp_2_addr = core_io_ptw_pmp_2_addr;
	assign ptw_io_dpath_pmp_2_mask = core_io_ptw_pmp_2_mask;
	assign ptw_io_dpath_pmp_3_cfg_l = core_io_ptw_pmp_3_cfg_l;
	assign ptw_io_dpath_pmp_3_cfg_a = core_io_ptw_pmp_3_cfg_a;
	assign ptw_io_dpath_pmp_3_cfg_x = core_io_ptw_pmp_3_cfg_x;
	assign ptw_io_dpath_pmp_3_cfg_w = core_io_ptw_pmp_3_cfg_w;
	assign ptw_io_dpath_pmp_3_cfg_r = core_io_ptw_pmp_3_cfg_r;
	assign ptw_io_dpath_pmp_3_addr = core_io_ptw_pmp_3_addr;
	assign ptw_io_dpath_pmp_3_mask = core_io_ptw_pmp_3_mask;
	assign ptw_io_dpath_pmp_4_cfg_l = core_io_ptw_pmp_4_cfg_l;
	assign ptw_io_dpath_pmp_4_cfg_a = core_io_ptw_pmp_4_cfg_a;
	assign ptw_io_dpath_pmp_4_cfg_x = core_io_ptw_pmp_4_cfg_x;
	assign ptw_io_dpath_pmp_4_cfg_w = core_io_ptw_pmp_4_cfg_w;
	assign ptw_io_dpath_pmp_4_cfg_r = core_io_ptw_pmp_4_cfg_r;
	assign ptw_io_dpath_pmp_4_addr = core_io_ptw_pmp_4_addr;
	assign ptw_io_dpath_pmp_4_mask = core_io_ptw_pmp_4_mask;
	assign ptw_io_dpath_pmp_5_cfg_l = core_io_ptw_pmp_5_cfg_l;
	assign ptw_io_dpath_pmp_5_cfg_a = core_io_ptw_pmp_5_cfg_a;
	assign ptw_io_dpath_pmp_5_cfg_x = core_io_ptw_pmp_5_cfg_x;
	assign ptw_io_dpath_pmp_5_cfg_w = core_io_ptw_pmp_5_cfg_w;
	assign ptw_io_dpath_pmp_5_cfg_r = core_io_ptw_pmp_5_cfg_r;
	assign ptw_io_dpath_pmp_5_addr = core_io_ptw_pmp_5_addr;
	assign ptw_io_dpath_pmp_5_mask = core_io_ptw_pmp_5_mask;
	assign ptw_io_dpath_pmp_6_cfg_l = core_io_ptw_pmp_6_cfg_l;
	assign ptw_io_dpath_pmp_6_cfg_a = core_io_ptw_pmp_6_cfg_a;
	assign ptw_io_dpath_pmp_6_cfg_x = core_io_ptw_pmp_6_cfg_x;
	assign ptw_io_dpath_pmp_6_cfg_w = core_io_ptw_pmp_6_cfg_w;
	assign ptw_io_dpath_pmp_6_cfg_r = core_io_ptw_pmp_6_cfg_r;
	assign ptw_io_dpath_pmp_6_addr = core_io_ptw_pmp_6_addr;
	assign ptw_io_dpath_pmp_6_mask = core_io_ptw_pmp_6_mask;
	assign ptw_io_dpath_pmp_7_cfg_l = core_io_ptw_pmp_7_cfg_l;
	assign ptw_io_dpath_pmp_7_cfg_a = core_io_ptw_pmp_7_cfg_a;
	assign ptw_io_dpath_pmp_7_cfg_x = core_io_ptw_pmp_7_cfg_x;
	assign ptw_io_dpath_pmp_7_cfg_w = core_io_ptw_pmp_7_cfg_w;
	assign ptw_io_dpath_pmp_7_cfg_r = core_io_ptw_pmp_7_cfg_r;
	assign ptw_io_dpath_pmp_7_addr = core_io_ptw_pmp_7_addr;
	assign ptw_io_dpath_pmp_7_mask = core_io_ptw_pmp_7_mask;
	assign ptw_io_dpath_customCSRs_csrs_0_value = core_io_ptw_customCSRs_csrs_0_value;
	assign core_clock = clock;
	assign core_reset = reset;
	assign core_io_hartid = broadcast_auto_out_0;
	assign core_io_interrupts_debug = intXbar_auto_int_out_0;
	assign core_io_interrupts_mtip = intXbar_auto_int_out_2;
	assign core_io_interrupts_msip = intXbar_auto_int_out_1;
	assign core_io_interrupts_meip = intXbar_auto_int_out_3;
	assign core_io_imem_resp_valid = frontend_io_cpu_resp_valid;
	assign core_io_imem_resp_bits_pc = frontend_io_cpu_resp_bits_pc;
	assign core_io_imem_resp_bits_data = frontend_io_cpu_resp_bits_data;
	assign core_io_imem_resp_bits_xcpt_ae_inst = frontend_io_cpu_resp_bits_xcpt_ae_inst;
	assign core_io_imem_resp_bits_replay = frontend_io_cpu_resp_bits_replay;
	assign core_io_dmem_req_ready = dcacheArb_io_requestor_0_req_ready;
	assign core_io_dmem_s2_nack = dcacheArb_io_requestor_0_s2_nack;
	assign core_io_dmem_resp_valid = dcacheArb_io_requestor_0_resp_valid;
	assign core_io_dmem_resp_bits_tag = dcacheArb_io_requestor_0_resp_bits_tag;
	assign core_io_dmem_resp_bits_data = dcacheArb_io_requestor_0_resp_bits_data;
	assign core_io_dmem_resp_bits_replay = dcacheArb_io_requestor_0_resp_bits_replay;
	assign core_io_dmem_resp_bits_has_data = dcacheArb_io_requestor_0_resp_bits_has_data;
	assign core_io_dmem_resp_bits_data_word_bypass = dcacheArb_io_requestor_0_resp_bits_data_word_bypass;
	assign core_io_dmem_replay_next = dcacheArb_io_requestor_0_replay_next;
	assign core_io_dmem_s2_xcpt_ma_ld = dcacheArb_io_requestor_0_s2_xcpt_ma_ld;
	assign core_io_dmem_s2_xcpt_ma_st = dcacheArb_io_requestor_0_s2_xcpt_ma_st;
	assign core_io_dmem_s2_xcpt_pf_ld = dcacheArb_io_requestor_0_s2_xcpt_pf_ld;
	assign core_io_dmem_s2_xcpt_pf_st = dcacheArb_io_requestor_0_s2_xcpt_pf_st;
	assign core_io_dmem_s2_xcpt_ae_ld = dcacheArb_io_requestor_0_s2_xcpt_ae_ld;
	assign core_io_dmem_s2_xcpt_ae_st = dcacheArb_io_requestor_0_s2_xcpt_ae_st;
	assign core_io_dmem_ordered = dcacheArb_io_requestor_0_ordered;
	assign core_io_dmem_perf_grant = dcacheArb_io_requestor_0_perf_grant;
	always @(posedge clock)
		if (reset)
			bundleOut_0_0_REG <= 1'h0;
		else
			bundleOut_0_0_REG <= core_io_wfi;
endmodule
module TileResetDomain (
	auto_tile_slave_in_a_ready,
	auto_tile_slave_in_a_valid,
	auto_tile_slave_in_a_bits_opcode,
	auto_tile_slave_in_a_bits_param,
	auto_tile_slave_in_a_bits_size,
	auto_tile_slave_in_a_bits_source,
	auto_tile_slave_in_a_bits_address,
	auto_tile_slave_in_a_bits_mask,
	auto_tile_slave_in_a_bits_data,
	auto_tile_slave_in_d_ready,
	auto_tile_slave_in_d_valid,
	auto_tile_slave_in_d_bits_opcode,
	auto_tile_slave_in_d_bits_size,
	auto_tile_slave_in_d_bits_source,
	auto_tile_slave_in_d_bits_data,
	auto_tile_wfi_out_0,
	auto_tile_int_local_in_2_0,
	auto_tile_int_local_in_1_0,
	auto_tile_int_local_in_1_1,
	auto_tile_int_local_in_0_0,
	auto_tile_hartid_in,
	auto_tile_tl_other_masters_out_a_ready,
	auto_tile_tl_other_masters_out_a_valid,
	auto_tile_tl_other_masters_out_a_bits_opcode,
	auto_tile_tl_other_masters_out_a_bits_param,
	auto_tile_tl_other_masters_out_a_bits_size,
	auto_tile_tl_other_masters_out_a_bits_source,
	auto_tile_tl_other_masters_out_a_bits_address,
	auto_tile_tl_other_masters_out_a_bits_mask,
	auto_tile_tl_other_masters_out_a_bits_data,
	auto_tile_tl_other_masters_out_d_ready,
	auto_tile_tl_other_masters_out_d_valid,
	auto_tile_tl_other_masters_out_d_bits_opcode,
	auto_tile_tl_other_masters_out_d_bits_param,
	auto_tile_tl_other_masters_out_d_bits_size,
	auto_tile_tl_other_masters_out_d_bits_source,
	auto_tile_tl_other_masters_out_d_bits_sink,
	auto_tile_tl_other_masters_out_d_bits_denied,
	auto_tile_tl_other_masters_out_d_bits_data,
	auto_tile_tl_other_masters_out_d_bits_corrupt,
	auto_clock_in_clock,
	auto_clock_in_reset
);
	output wire auto_tile_slave_in_a_ready;
	input auto_tile_slave_in_a_valid;
	input [2:0] auto_tile_slave_in_a_bits_opcode;
	input [2:0] auto_tile_slave_in_a_bits_param;
	input [2:0] auto_tile_slave_in_a_bits_size;
	input [2:0] auto_tile_slave_in_a_bits_source;
	input [31:0] auto_tile_slave_in_a_bits_address;
	input [3:0] auto_tile_slave_in_a_bits_mask;
	input [31:0] auto_tile_slave_in_a_bits_data;
	input auto_tile_slave_in_d_ready;
	output wire auto_tile_slave_in_d_valid;
	output wire [2:0] auto_tile_slave_in_d_bits_opcode;
	output wire [2:0] auto_tile_slave_in_d_bits_size;
	output wire [2:0] auto_tile_slave_in_d_bits_source;
	output wire [31:0] auto_tile_slave_in_d_bits_data;
	output wire auto_tile_wfi_out_0;
	input auto_tile_int_local_in_2_0;
	input auto_tile_int_local_in_1_0;
	input auto_tile_int_local_in_1_1;
	input auto_tile_int_local_in_0_0;
	input auto_tile_hartid_in;
	input auto_tile_tl_other_masters_out_a_ready;
	output wire auto_tile_tl_other_masters_out_a_valid;
	output wire [2:0] auto_tile_tl_other_masters_out_a_bits_opcode;
	output wire [2:0] auto_tile_tl_other_masters_out_a_bits_param;
	output wire [3:0] auto_tile_tl_other_masters_out_a_bits_size;
	output wire auto_tile_tl_other_masters_out_a_bits_source;
	output wire [31:0] auto_tile_tl_other_masters_out_a_bits_address;
	output wire [3:0] auto_tile_tl_other_masters_out_a_bits_mask;
	output wire [31:0] auto_tile_tl_other_masters_out_a_bits_data;
	output wire auto_tile_tl_other_masters_out_d_ready;
	input auto_tile_tl_other_masters_out_d_valid;
	input [2:0] auto_tile_tl_other_masters_out_d_bits_opcode;
	input [1:0] auto_tile_tl_other_masters_out_d_bits_param;
	input [3:0] auto_tile_tl_other_masters_out_d_bits_size;
	input auto_tile_tl_other_masters_out_d_bits_source;
	input auto_tile_tl_other_masters_out_d_bits_sink;
	input auto_tile_tl_other_masters_out_d_bits_denied;
	input [31:0] auto_tile_tl_other_masters_out_d_bits_data;
	input auto_tile_tl_other_masters_out_d_bits_corrupt;
	input auto_clock_in_clock;
	input auto_clock_in_reset;
	wire tile_clock;
	wire tile_reset;
	wire tile_auto_slave_in_a_ready;
	wire tile_auto_slave_in_a_valid;
	wire [2:0] tile_auto_slave_in_a_bits_opcode;
	wire [2:0] tile_auto_slave_in_a_bits_param;
	wire [2:0] tile_auto_slave_in_a_bits_size;
	wire [2:0] tile_auto_slave_in_a_bits_source;
	wire [31:0] tile_auto_slave_in_a_bits_address;
	wire [3:0] tile_auto_slave_in_a_bits_mask;
	wire [31:0] tile_auto_slave_in_a_bits_data;
	wire tile_auto_slave_in_d_ready;
	wire tile_auto_slave_in_d_valid;
	wire [2:0] tile_auto_slave_in_d_bits_opcode;
	wire [2:0] tile_auto_slave_in_d_bits_size;
	wire [2:0] tile_auto_slave_in_d_bits_source;
	wire [31:0] tile_auto_slave_in_d_bits_data;
	wire tile_auto_wfi_out_0;
	wire tile_auto_int_local_in_2_0;
	wire tile_auto_int_local_in_1_0;
	wire tile_auto_int_local_in_1_1;
	wire tile_auto_int_local_in_0_0;
	wire tile_auto_hartid_in;
	wire tile_auto_tl_other_masters_out_a_ready;
	wire tile_auto_tl_other_masters_out_a_valid;
	wire [2:0] tile_auto_tl_other_masters_out_a_bits_opcode;
	wire [2:0] tile_auto_tl_other_masters_out_a_bits_param;
	wire [3:0] tile_auto_tl_other_masters_out_a_bits_size;
	wire tile_auto_tl_other_masters_out_a_bits_source;
	wire [31:0] tile_auto_tl_other_masters_out_a_bits_address;
	wire [3:0] tile_auto_tl_other_masters_out_a_bits_mask;
	wire [31:0] tile_auto_tl_other_masters_out_a_bits_data;
	wire tile_auto_tl_other_masters_out_d_ready;
	wire tile_auto_tl_other_masters_out_d_valid;
	wire [2:0] tile_auto_tl_other_masters_out_d_bits_opcode;
	wire [1:0] tile_auto_tl_other_masters_out_d_bits_param;
	wire [3:0] tile_auto_tl_other_masters_out_d_bits_size;
	wire tile_auto_tl_other_masters_out_d_bits_source;
	wire tile_auto_tl_other_masters_out_d_bits_sink;
	wire tile_auto_tl_other_masters_out_d_bits_denied;
	wire [31:0] tile_auto_tl_other_masters_out_d_bits_data;
	wire tile_auto_tl_other_masters_out_d_bits_corrupt;
	RocketTile tile(
		.clock(tile_clock),
		.reset(tile_reset),
		.auto_slave_in_a_ready(tile_auto_slave_in_a_ready),
		.auto_slave_in_a_valid(tile_auto_slave_in_a_valid),
		.auto_slave_in_a_bits_opcode(tile_auto_slave_in_a_bits_opcode),
		.auto_slave_in_a_bits_param(tile_auto_slave_in_a_bits_param),
		.auto_slave_in_a_bits_size(tile_auto_slave_in_a_bits_size),
		.auto_slave_in_a_bits_source(tile_auto_slave_in_a_bits_source),
		.auto_slave_in_a_bits_address(tile_auto_slave_in_a_bits_address),
		.auto_slave_in_a_bits_mask(tile_auto_slave_in_a_bits_mask),
		.auto_slave_in_a_bits_data(tile_auto_slave_in_a_bits_data),
		.auto_slave_in_d_ready(tile_auto_slave_in_d_ready),
		.auto_slave_in_d_valid(tile_auto_slave_in_d_valid),
		.auto_slave_in_d_bits_opcode(tile_auto_slave_in_d_bits_opcode),
		.auto_slave_in_d_bits_size(tile_auto_slave_in_d_bits_size),
		.auto_slave_in_d_bits_source(tile_auto_slave_in_d_bits_source),
		.auto_slave_in_d_bits_data(tile_auto_slave_in_d_bits_data),
		.auto_wfi_out_0(tile_auto_wfi_out_0),
		.auto_int_local_in_2_0(tile_auto_int_local_in_2_0),
		.auto_int_local_in_1_0(tile_auto_int_local_in_1_0),
		.auto_int_local_in_1_1(tile_auto_int_local_in_1_1),
		.auto_int_local_in_0_0(tile_auto_int_local_in_0_0),
		.auto_hartid_in(tile_auto_hartid_in),
		.auto_tl_other_masters_out_a_ready(tile_auto_tl_other_masters_out_a_ready),
		.auto_tl_other_masters_out_a_valid(tile_auto_tl_other_masters_out_a_valid),
		.auto_tl_other_masters_out_a_bits_opcode(tile_auto_tl_other_masters_out_a_bits_opcode),
		.auto_tl_other_masters_out_a_bits_param(tile_auto_tl_other_masters_out_a_bits_param),
		.auto_tl_other_masters_out_a_bits_size(tile_auto_tl_other_masters_out_a_bits_size),
		.auto_tl_other_masters_out_a_bits_source(tile_auto_tl_other_masters_out_a_bits_source),
		.auto_tl_other_masters_out_a_bits_address(tile_auto_tl_other_masters_out_a_bits_address),
		.auto_tl_other_masters_out_a_bits_mask(tile_auto_tl_other_masters_out_a_bits_mask),
		.auto_tl_other_masters_out_a_bits_data(tile_auto_tl_other_masters_out_a_bits_data),
		.auto_tl_other_masters_out_d_ready(tile_auto_tl_other_masters_out_d_ready),
		.auto_tl_other_masters_out_d_valid(tile_auto_tl_other_masters_out_d_valid),
		.auto_tl_other_masters_out_d_bits_opcode(tile_auto_tl_other_masters_out_d_bits_opcode),
		.auto_tl_other_masters_out_d_bits_param(tile_auto_tl_other_masters_out_d_bits_param),
		.auto_tl_other_masters_out_d_bits_size(tile_auto_tl_other_masters_out_d_bits_size),
		.auto_tl_other_masters_out_d_bits_source(tile_auto_tl_other_masters_out_d_bits_source),
		.auto_tl_other_masters_out_d_bits_sink(tile_auto_tl_other_masters_out_d_bits_sink),
		.auto_tl_other_masters_out_d_bits_denied(tile_auto_tl_other_masters_out_d_bits_denied),
		.auto_tl_other_masters_out_d_bits_data(tile_auto_tl_other_masters_out_d_bits_data),
		.auto_tl_other_masters_out_d_bits_corrupt(tile_auto_tl_other_masters_out_d_bits_corrupt)
	);
	assign auto_tile_slave_in_a_ready = tile_auto_slave_in_a_ready;
	assign auto_tile_slave_in_d_valid = tile_auto_slave_in_d_valid;
	assign auto_tile_slave_in_d_bits_opcode = tile_auto_slave_in_d_bits_opcode;
	assign auto_tile_slave_in_d_bits_size = tile_auto_slave_in_d_bits_size;
	assign auto_tile_slave_in_d_bits_source = tile_auto_slave_in_d_bits_source;
	assign auto_tile_slave_in_d_bits_data = tile_auto_slave_in_d_bits_data;
	assign auto_tile_wfi_out_0 = tile_auto_wfi_out_0;
	assign auto_tile_tl_other_masters_out_a_valid = tile_auto_tl_other_masters_out_a_valid;
	assign auto_tile_tl_other_masters_out_a_bits_opcode = tile_auto_tl_other_masters_out_a_bits_opcode;
	assign auto_tile_tl_other_masters_out_a_bits_param = tile_auto_tl_other_masters_out_a_bits_param;
	assign auto_tile_tl_other_masters_out_a_bits_size = tile_auto_tl_other_masters_out_a_bits_size;
	assign auto_tile_tl_other_masters_out_a_bits_source = tile_auto_tl_other_masters_out_a_bits_source;
	assign auto_tile_tl_other_masters_out_a_bits_address = tile_auto_tl_other_masters_out_a_bits_address;
	assign auto_tile_tl_other_masters_out_a_bits_mask = tile_auto_tl_other_masters_out_a_bits_mask;
	assign auto_tile_tl_other_masters_out_a_bits_data = tile_auto_tl_other_masters_out_a_bits_data;
	assign auto_tile_tl_other_masters_out_d_ready = tile_auto_tl_other_masters_out_d_ready;
	assign tile_clock = auto_clock_in_clock;
	assign tile_reset = auto_clock_in_reset;
	assign tile_auto_slave_in_a_valid = auto_tile_slave_in_a_valid;
	assign tile_auto_slave_in_a_bits_opcode = auto_tile_slave_in_a_bits_opcode;
	assign tile_auto_slave_in_a_bits_param = auto_tile_slave_in_a_bits_param;
	assign tile_auto_slave_in_a_bits_size = auto_tile_slave_in_a_bits_size;
	assign tile_auto_slave_in_a_bits_source = auto_tile_slave_in_a_bits_source;
	assign tile_auto_slave_in_a_bits_address = auto_tile_slave_in_a_bits_address;
	assign tile_auto_slave_in_a_bits_mask = auto_tile_slave_in_a_bits_mask;
	assign tile_auto_slave_in_a_bits_data = auto_tile_slave_in_a_bits_data;
	assign tile_auto_slave_in_d_ready = auto_tile_slave_in_d_ready;
	assign tile_auto_int_local_in_2_0 = auto_tile_int_local_in_2_0;
	assign tile_auto_int_local_in_1_0 = auto_tile_int_local_in_1_0;
	assign tile_auto_int_local_in_1_1 = auto_tile_int_local_in_1_1;
	assign tile_auto_int_local_in_0_0 = auto_tile_int_local_in_0_0;
	assign tile_auto_hartid_in = auto_tile_hartid_in;
	assign tile_auto_tl_other_masters_out_a_ready = auto_tile_tl_other_masters_out_a_ready;
	assign tile_auto_tl_other_masters_out_d_valid = auto_tile_tl_other_masters_out_d_valid;
	assign tile_auto_tl_other_masters_out_d_bits_opcode = auto_tile_tl_other_masters_out_d_bits_opcode;
	assign tile_auto_tl_other_masters_out_d_bits_param = auto_tile_tl_other_masters_out_d_bits_param;
	assign tile_auto_tl_other_masters_out_d_bits_size = auto_tile_tl_other_masters_out_d_bits_size;
	assign tile_auto_tl_other_masters_out_d_bits_source = auto_tile_tl_other_masters_out_d_bits_source;
	assign tile_auto_tl_other_masters_out_d_bits_sink = auto_tile_tl_other_masters_out_d_bits_sink;
	assign tile_auto_tl_other_masters_out_d_bits_denied = auto_tile_tl_other_masters_out_d_bits_denied;
	assign tile_auto_tl_other_masters_out_d_bits_data = auto_tile_tl_other_masters_out_d_bits_data;
	assign tile_auto_tl_other_masters_out_d_bits_corrupt = auto_tile_tl_other_masters_out_d_bits_corrupt;
endmodule
module FixedClockBroadcast_4 (
	auto_in_clock,
	auto_in_reset,
	auto_out_clock,
	auto_out_reset
);
	input auto_in_clock;
	input auto_in_reset;
	output wire auto_out_clock;
	output wire auto_out_reset;
	assign auto_out_clock = auto_in_clock;
	assign auto_out_reset = auto_in_reset;
endmodule
module TLBuffer_13 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_param = auto_out_d_bits_param;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_sink = auto_out_d_bits_sink;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module TLMonitor_33 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [3:0] io_in_a_bits_size;
	input io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_1 = ~io_in_a_bits_source;
	wire source_ok = io_in_a_bits_source | _source_ok_T_1;
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << io_in_a_bits_size;
	wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0];
	wire [31:0] _GEN_71 = {20'd0, is_aligned_mask};
	wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 32'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 4'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire [32:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_24 = io_in_a_bits_opcode == 3'h6;
	wire _T_26 = io_in_a_bits_size <= 4'hc;
	wire _T_31 = _T_26 & source_ok;
	wire [32:0] _T_37 = $signed(_T_7) & -33'sh000005000;
	wire _T_38 = $signed(_T_37) == 33'sh000000000;
	wire [31:0] _T_39 = io_in_a_bits_address ^ 32'h00003000;
	wire [32:0] _T_40 = {1'b0, $signed(_T_39)};
	wire [32:0] _T_42 = $signed(_T_40) & -33'sh000001000;
	wire _T_43 = $signed(_T_42) == 33'sh000000000;
	wire [31:0] _T_44 = io_in_a_bits_address ^ 32'h00010000;
	wire [32:0] _T_45 = {1'b0, $signed(_T_44)};
	wire [32:0] _T_47 = $signed(_T_45) & -33'sh000010000;
	wire _T_48 = $signed(_T_47) == 33'sh000000000;
	wire [31:0] _T_49 = io_in_a_bits_address ^ 32'h00020000;
	wire [32:0] _T_50 = {1'b0, $signed(_T_49)};
	wire [32:0] _T_52 = $signed(_T_50) & -33'sh000010000;
	wire _T_53 = $signed(_T_52) == 33'sh000000000;
	wire [31:0] _T_54 = io_in_a_bits_address ^ 32'h00100000;
	wire [32:0] _T_55 = {1'b0, $signed(_T_54)};
	wire [32:0] _T_57 = $signed(_T_55) & -33'sh000011000;
	wire _T_58 = $signed(_T_57) == 33'sh000000000;
	wire [31:0] _T_59 = io_in_a_bits_address ^ 32'h02000000;
	wire [32:0] _T_60 = {1'b0, $signed(_T_59)};
	wire [32:0] _T_62 = $signed(_T_60) & -33'sh000010000;
	wire _T_63 = $signed(_T_62) == 33'sh000000000;
	wire [31:0] _T_64 = io_in_a_bits_address ^ 32'h0c000000;
	wire [32:0] _T_65 = {1'b0, $signed(_T_64)};
	wire [32:0] _T_67 = $signed(_T_65) & -33'sh004000000;
	wire _T_68 = $signed(_T_67) == 33'sh000000000;
	wire [31:0] _T_69 = io_in_a_bits_address ^ 32'h10000000;
	wire [32:0] _T_70 = {1'b0, $signed(_T_69)};
	wire [32:0] _T_72 = $signed(_T_70) & -33'sh000001000;
	wire _T_73 = $signed(_T_72) == 33'sh000000000;
	wire [31:0] _T_74 = io_in_a_bits_address ^ 32'h54000000;
	wire [32:0] _T_75 = {1'b0, $signed(_T_74)};
	wire [32:0] _T_77 = $signed(_T_75) & -33'sh000001000;
	wire _T_78 = $signed(_T_77) == 33'sh000000000;
	wire [31:0] _T_79 = io_in_a_bits_address ^ 32'h80000000;
	wire [32:0] _T_80 = {1'b0, $signed(_T_79)};
	wire [32:0] _T_82 = $signed(_T_80) & -33'sh000004000;
	wire _T_83 = $signed(_T_82) == 33'sh000000000;
	wire _T_178 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_182 = ~io_in_a_bits_mask;
	wire _T_183 = _T_182 == 4'h0;
	wire _T_191 = io_in_a_bits_opcode == 3'h7;
	wire _T_349 = io_in_a_bits_param != 3'h0;
	wire _T_362 = io_in_a_bits_opcode == 3'h4;
	wire _T_383 = _T_26 & _T_43;
	wire _T_385 = io_in_a_bits_size <= 4'h6;
	wire _T_440 = (((((((_T_38 | _T_48) | _T_53) | _T_58) | _T_63) | _T_68) | _T_73) | _T_78) | _T_83;
	wire _T_441 = _T_385 & _T_440;
	wire _T_443 = _T_383 | _T_441;
	wire _T_453 = io_in_a_bits_param == 3'h0;
	wire _T_457 = io_in_a_bits_mask == mask;
	wire _T_465 = io_in_a_bits_opcode == 3'h0;
	wire _T_528 = (((((_T_38 | _T_58) | _T_63) | _T_68) | _T_73) | _T_78) | _T_83;
	wire _T_529 = _T_385 & _T_528;
	wire _T_544 = _T_383 | _T_529;
	wire _T_546 = _T_31 & _T_544;
	wire _T_564 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_659 = ~mask;
	wire [3:0] _T_660 = io_in_a_bits_mask & _T_659;
	wire _T_661 = _T_660 == 4'h0;
	wire _T_665 = io_in_a_bits_opcode == 3'h2;
	wire _T_675 = io_in_a_bits_size <= 4'h2;
	wire _T_724 = ((((((_T_38 | _T_43) | _T_58) | _T_63) | _T_68) | _T_73) | _T_78) | _T_83;
	wire _T_725 = _T_675 & _T_724;
	wire _T_741 = _T_31 & _T_725;
	wire _T_751 = io_in_a_bits_param <= 3'h4;
	wire _T_759 = io_in_a_bits_opcode == 3'h3;
	wire _T_845 = io_in_a_bits_param <= 3'h3;
	wire _T_853 = io_in_a_bits_opcode == 3'h5;
	wire _T_929 = _T_31 & _T_383;
	wire _T_939 = io_in_a_bits_param <= 3'h1;
	wire _T_951 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_3 = ~io_in_d_bits_source;
	wire source_ok_1 = io_in_d_bits_source | _source_ok_T_3;
	wire _T_955 = io_in_d_bits_opcode == 3'h6;
	wire _T_959 = io_in_d_bits_size >= 4'h2;
	wire _T_963 = io_in_d_bits_param == 2'h0;
	wire _T_967 = ~io_in_d_bits_corrupt;
	wire _T_971 = ~io_in_d_bits_denied;
	wire _T_975 = io_in_d_bits_opcode == 3'h4;
	wire _T_986 = io_in_d_bits_param <= 2'h2;
	wire _T_990 = io_in_d_bits_param != 2'h2;
	wire _T_1003 = io_in_d_bits_opcode == 3'h5;
	wire _T_1023 = _T_971 | io_in_d_bits_corrupt;
	wire _T_1032 = io_in_d_bits_opcode == 3'h0;
	wire _T_1049 = io_in_d_bits_opcode == 3'h1;
	wire _T_1067 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [9:0] a_first_counter;
	wire [9:0] a_first_counter1 = a_first_counter - 10'h001;
	wire a_first = a_first_counter == 10'h000;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [3:0] size;
	reg source;
	reg [31:0] address;
	wire _T_1097 = io_in_a_valid & ~a_first;
	wire _T_1098 = io_in_a_bits_opcode == opcode;
	wire _T_1102 = io_in_a_bits_param == param;
	wire _T_1106 = io_in_a_bits_size == size;
	wire _T_1110 = io_in_a_bits_source == source;
	wire _T_1114 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << io_in_d_bits_size;
	wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0];
	wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [9:0] d_first_counter;
	wire [9:0] d_first_counter1 = d_first_counter - 10'h001;
	wire d_first = d_first_counter == 10'h000;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg source_1;
	reg sink;
	reg denied;
	wire _T_1121 = io_in_d_valid & ~d_first;
	wire _T_1122 = io_in_d_bits_opcode == opcode_1;
	wire _T_1126 = io_in_d_bits_param == param_1;
	wire _T_1130 = io_in_d_bits_size == size_1;
	wire _T_1134 = io_in_d_bits_source == source_1;
	wire _T_1138 = io_in_d_bits_sink == sink;
	wire _T_1142 = io_in_d_bits_denied == denied;
	reg [1:0] inflight;
	reg [7:0] inflight_opcodes;
	reg [15:0] inflight_sizes;
	reg [9:0] a_first_counter_1;
	wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h001;
	wire a_first_1 = a_first_counter_1 == 10'h000;
	reg [9:0] d_first_counter_1;
	wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h001;
	wire d_first_1 = d_first_counter_1 == 10'h000;
	wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [3:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [7:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_73 = {8'd0, _a_opcode_lookup_T_1};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0};
	wire [15:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T;
	wire [15:0] _a_size_lookup_T_5 = 16'h0100 - 16'h0001;
	wire [15:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _a_size_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_1148 = io_in_a_valid & a_first_1;
	wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source;
	wire [1:0] a_set_wo_ready = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire _T_1151 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h01;
	wire [2:0] _GEN_76 = {io_in_a_bits_source, 2'h0};
	wire [3:0] _a_opcodes_set_T = {1'd0, _GEN_76};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _GEN_1 = {15'd0, a_opcodes_set_interm};
	wire [18:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0};
	wire [4:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h00);
	wire [19:0] _GEN_2 = {15'd0, a_sizes_set_interm};
	wire [19:0] _a_sizes_set_T_1 = _GEN_2 << _a_sizes_set_T;
	wire [1:0] _T_1153 = inflight >> io_in_a_bits_source;
	wire _T_1155 = ~_T_1153[0];
	wire [1:0] a_set = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire [18:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [19:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 20'h00000);
	wire _T_1159 = io_in_d_valid & d_first_1;
	wire _T_1161 = ~_T_955;
	wire _T_1162 = (io_in_d_valid & d_first_1) & ~_T_955;
	wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source;
	wire [1:0] d_clr_wo_ready = ((io_in_d_valid & d_first_1) & ~_T_955 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_3 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [30:0] _GEN_4 = {15'd0, _a_size_lookup_T_5};
	wire [30:0] _d_sizes_clr_T_5 = _GEN_4 << _a_size_lookup_T;
	wire [1:0] d_clr = ((_d_first_T & d_first_1) & _T_1161 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_1161 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [30:0] _GEN_24 = ((_d_first_T & d_first_1) & _T_1161 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_1148 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [1:0] _T_1172 = inflight >> io_in_d_bits_source;
	wire _T_1174 = _T_1172[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_1179 = io_in_d_bits_opcode == _GEN_40;
	wire _T_1180 = (io_in_d_bits_opcode == _GEN_32) | _T_1179;
	wire _T_1184 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_1191 = io_in_d_bits_opcode == _GEN_56;
	wire _T_1192 = (io_in_d_bits_opcode == _GEN_48) | _T_1191;
	wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
	wire [7:0] _GEN_78 = {4'd0, io_in_d_bits_size};
	wire _T_1196 = _GEN_78 == a_size_lookup;
	wire _T_1206 = (((_T_1159 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_1161;
	wire _T_1208 = ~io_in_d_ready | io_in_a_ready;
	wire _T_1215 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [1:0] _inflight_T = inflight | a_set;
	wire [1:0] _inflight_T_1 = ~d_clr;
	wire [1:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [7:0] a_opcodes_set = _GEN_19[7:0];
	wire [7:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [7:0] d_opcodes_clr = _GEN_23[7:0];
	wire [7:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [7:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [15:0] a_sizes_set = _GEN_20[15:0];
	wire [15:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [15:0] d_sizes_clr = _GEN_24[15:0];
	wire [15:0] _inflight_sizes_T_1 = ~d_sizes_clr;
	wire [15:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1;
	reg [31:0] watchdog;
	wire _T_1224 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [1:0] inflight_1;
	reg [15:0] inflight_sizes_1;
	reg [9:0] d_first_counter_2;
	wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h001;
	wire d_first_2 = d_first_counter_2 == 10'h000;
	wire [15:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T;
	wire [15:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _a_size_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_1250 = (io_in_d_valid & d_first_2) & _T_955;
	wire [1:0] d_clr_1 = ((_d_first_T & d_first_2) & _T_955 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_69 = ((_d_first_T & d_first_2) & _T_955 ? _d_sizes_clr_T_5 : 31'h00000000);
	wire [1:0] _T_1258 = inflight_1 >> io_in_d_bits_source;
	wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
	wire _T_1268 = _GEN_78 == c_size_lookup;
	wire [1:0] _inflight_T_4 = ~d_clr_1;
	wire [1:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [15:0] d_sizes_clr_1 = _GEN_69[15:0];
	wire [15:0] _inflight_sizes_T_4 = ~d_sizes_clr_1;
	wire [15:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4;
	reg [31:0] watchdog_1;
	wire _T_1293 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 10'h000;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 10'h000;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 10'h000;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 10'h000;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 2'h0;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 8'h00;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 16'h0000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 10'h000;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 10'h000;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 10'h000;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 10'h000;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 2'h0;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 16'h0000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 10'h000;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 10'h000;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLBuffer_14 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [3:0] auto_in_a_bits_size;
	input auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [3:0] monitor_io_in_a_bits_size;
	wire monitor_io_in_a_bits_source;
	wire [31:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [3:0] monitor_io_in_d_bits_size;
	wire monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire bundleOut_0_a_q_clock;
	wire bundleOut_0_a_q_reset;
	wire bundleOut_0_a_q_io_enq_ready;
	wire bundleOut_0_a_q_io_enq_valid;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_param;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_size;
	wire bundleOut_0_a_q_io_enq_bits_source;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_data;
	wire bundleOut_0_a_q_io_enq_bits_corrupt;
	wire bundleOut_0_a_q_io_deq_ready;
	wire bundleOut_0_a_q_io_deq_valid;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_param;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_size;
	wire bundleOut_0_a_q_io_deq_bits_source;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_data;
	wire bundleOut_0_a_q_io_deq_bits_corrupt;
	wire bundleIn_0_d_q_clock;
	wire bundleIn_0_d_q_reset;
	wire bundleIn_0_d_q_io_enq_ready;
	wire bundleIn_0_d_q_io_enq_valid;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_enq_bits_param;
	wire [3:0] bundleIn_0_d_q_io_enq_bits_size;
	wire bundleIn_0_d_q_io_enq_bits_source;
	wire bundleIn_0_d_q_io_enq_bits_sink;
	wire bundleIn_0_d_q_io_enq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_enq_bits_data;
	wire bundleIn_0_d_q_io_enq_bits_corrupt;
	wire bundleIn_0_d_q_io_deq_ready;
	wire bundleIn_0_d_q_io_deq_valid;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_param;
	wire [3:0] bundleIn_0_d_q_io_deq_bits_size;
	wire bundleIn_0_d_q_io_deq_bits_source;
	wire bundleIn_0_d_q_io_deq_bits_sink;
	wire bundleIn_0_d_q_io_deq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_deq_bits_data;
	wire bundleIn_0_d_q_io_deq_bits_corrupt;
	TLMonitor_33 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Queue_4 bundleOut_0_a_q(
		.clock(bundleOut_0_a_q_clock),
		.reset(bundleOut_0_a_q_reset),
		.io_enq_ready(bundleOut_0_a_q_io_enq_ready),
		.io_enq_valid(bundleOut_0_a_q_io_enq_valid),
		.io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
		.io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
		.io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
		.io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
		.io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
		.io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleOut_0_a_q_io_deq_ready),
		.io_deq_valid(bundleOut_0_a_q_io_deq_valid),
		.io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
		.io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
		.io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
		.io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
		.io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
		.io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
	);
	Queue_5 bundleIn_0_d_q(
		.clock(bundleIn_0_d_q_clock),
		.reset(bundleIn_0_d_q_reset),
		.io_enq_ready(bundleIn_0_d_q_io_enq_ready),
		.io_enq_valid(bundleIn_0_d_q_io_enq_valid),
		.io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
		.io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
		.io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
		.io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
		.io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
		.io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleIn_0_d_q_io_deq_ready),
		.io_deq_valid(bundleIn_0_d_q_io_deq_valid),
		.io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
		.io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
		.io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
		.io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
		.io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
		.io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data;
	assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid;
	assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode;
	assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param;
	assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size;
	assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source;
	assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address;
	assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask;
	assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data;
	assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt;
	assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign bundleOut_0_a_q_clock = clock;
	assign bundleOut_0_a_q_reset = reset;
	assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid;
	assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param;
	assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size;
	assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source;
	assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address;
	assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask;
	assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data;
	assign bundleOut_0_a_q_io_enq_bits_corrupt = 1'h0;
	assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready;
	assign bundleIn_0_d_q_clock = clock;
	assign bundleIn_0_d_q_reset = reset;
	assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid;
	assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign bundleIn_0_d_q_io_enq_bits_param = auto_out_d_bits_param;
	assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size;
	assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source;
	assign bundleIn_0_d_q_io_enq_bits_sink = auto_out_d_bits_sink;
	assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied;
	assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data;
	assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt;
	assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready;
endmodule
module TLBuffer_15 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module Queue_19 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_data,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_data
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [31:0] io_enq_bits_address;
	input [3:0] io_enq_bits_mask;
	input [31:0] io_enq_bits_data;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [31:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire [31:0] io_deq_bits_data;
	reg [2:0] ram_opcode [0:1];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [2:0] ram_param [0:1];
	wire ram_param_io_deq_bits_MPORT_en;
	wire ram_param_io_deq_bits_MPORT_addr;
	wire [2:0] ram_param_io_deq_bits_MPORT_data;
	wire [2:0] ram_param_MPORT_data;
	wire ram_param_MPORT_addr;
	wire ram_param_MPORT_mask;
	wire ram_param_MPORT_en;
	reg [2:0] ram_size [0:1];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [2:0] ram_size_io_deq_bits_MPORT_data;
	wire [2:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg [2:0] ram_source [0:1];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire [2:0] ram_source_io_deq_bits_MPORT_data;
	wire [2:0] ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg [31:0] ram_address [0:1];
	wire ram_address_io_deq_bits_MPORT_en;
	wire ram_address_io_deq_bits_MPORT_addr;
	wire [31:0] ram_address_io_deq_bits_MPORT_data;
	wire [31:0] ram_address_MPORT_data;
	wire ram_address_MPORT_addr;
	wire ram_address_MPORT_mask;
	wire ram_address_MPORT_en;
	reg [3:0] ram_mask [0:1];
	wire ram_mask_io_deq_bits_MPORT_en;
	wire ram_mask_io_deq_bits_MPORT_addr;
	wire [3:0] ram_mask_io_deq_bits_MPORT_data;
	wire [3:0] ram_mask_MPORT_data;
	wire ram_mask_MPORT_addr;
	wire ram_mask_MPORT_mask;
	wire ram_mask_MPORT_en;
	reg [31:0] ram_data [0:1];
	wire ram_data_io_deq_bits_MPORT_en;
	wire ram_data_io_deq_bits_MPORT_addr;
	wire [31:0] ram_data_io_deq_bits_MPORT_data;
	wire [31:0] ram_data_MPORT_data;
	wire ram_data_MPORT_addr;
	wire ram_data_MPORT_mask;
	wire ram_data_MPORT_en;
	reg value;
	reg value_1;
	reg maybe_full;
	wire ptr_match = value == value_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = value;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_param_io_deq_bits_MPORT_en = 1'h1;
	assign ram_param_io_deq_bits_MPORT_addr = value_1;
	assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr];
	assign ram_param_MPORT_data = io_enq_bits_param;
	assign ram_param_MPORT_addr = value;
	assign ram_param_MPORT_mask = 1'h1;
	assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = value_1;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = value;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = value_1;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = value;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_address_io_deq_bits_MPORT_en = 1'h1;
	assign ram_address_io_deq_bits_MPORT_addr = value_1;
	assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr];
	assign ram_address_MPORT_data = io_enq_bits_address;
	assign ram_address_MPORT_addr = value;
	assign ram_address_MPORT_mask = 1'h1;
	assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
	assign ram_mask_io_deq_bits_MPORT_addr = value_1;
	assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr];
	assign ram_mask_MPORT_data = io_enq_bits_mask;
	assign ram_mask_MPORT_addr = value;
	assign ram_mask_MPORT_mask = 1'h1;
	assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_data_io_deq_bits_MPORT_en = 1'h1;
	assign ram_data_io_deq_bits_MPORT_addr = value_1;
	assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr];
	assign ram_data_MPORT_data = io_enq_bits_data;
	assign ram_data_MPORT_addr = value;
	assign ram_data_MPORT_mask = 1'h1;
	assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data;
	assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data;
	assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_param_MPORT_en & ram_param_MPORT_mask)
			ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (ram_address_MPORT_en & ram_address_MPORT_mask)
			ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data;
		if (ram_mask_MPORT_en & ram_mask_MPORT_mask)
			ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data;
		if (ram_data_MPORT_en & ram_data_MPORT_mask)
			ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data;
		if (reset)
			value <= 1'h0;
		else if (do_enq)
			value <= value + 1'h1;
		if (reset)
			value_1 <= 1'h0;
		else if (do_deq)
			value_1 <= value_1 + 1'h1;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module TLBuffer_16 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	wire bundleOut_0_a_q_clock;
	wire bundleOut_0_a_q_reset;
	wire bundleOut_0_a_q_io_enq_ready;
	wire bundleOut_0_a_q_io_enq_valid;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_param;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_size;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_source;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_enq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_enq_bits_data;
	wire bundleOut_0_a_q_io_deq_ready;
	wire bundleOut_0_a_q_io_deq_valid;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_param;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_size;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_source;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_address;
	wire [3:0] bundleOut_0_a_q_io_deq_bits_mask;
	wire [31:0] bundleOut_0_a_q_io_deq_bits_data;
	wire bundleIn_0_d_q_clock;
	wire bundleIn_0_d_q_reset;
	wire bundleIn_0_d_q_io_enq_ready;
	wire bundleIn_0_d_q_io_enq_valid;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_enq_bits_param;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_size;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_source;
	wire bundleIn_0_d_q_io_enq_bits_sink;
	wire bundleIn_0_d_q_io_enq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_enq_bits_data;
	wire bundleIn_0_d_q_io_enq_bits_corrupt;
	wire bundleIn_0_d_q_io_deq_ready;
	wire bundleIn_0_d_q_io_deq_valid;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_param;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_size;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_source;
	wire bundleIn_0_d_q_io_deq_bits_sink;
	wire bundleIn_0_d_q_io_deq_bits_denied;
	wire [31:0] bundleIn_0_d_q_io_deq_bits_data;
	wire bundleIn_0_d_q_io_deq_bits_corrupt;
	Queue_19 bundleOut_0_a_q(
		.clock(bundleOut_0_a_q_clock),
		.reset(bundleOut_0_a_q_reset),
		.io_enq_ready(bundleOut_0_a_q_io_enq_ready),
		.io_enq_valid(bundleOut_0_a_q_io_enq_valid),
		.io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
		.io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
		.io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
		.io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
		.io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
		.io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
		.io_deq_ready(bundleOut_0_a_q_io_deq_ready),
		.io_deq_valid(bundleOut_0_a_q_io_deq_valid),
		.io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
		.io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
		.io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
		.io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
		.io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
		.io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data)
	);
	Queue_1 bundleIn_0_d_q(
		.clock(bundleIn_0_d_q_clock),
		.reset(bundleIn_0_d_q_reset),
		.io_enq_ready(bundleIn_0_d_q_io_enq_ready),
		.io_enq_valid(bundleIn_0_d_q_io_enq_valid),
		.io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
		.io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
		.io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
		.io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
		.io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
		.io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleIn_0_d_q_io_deq_ready),
		.io_deq_valid(bundleIn_0_d_q_io_deq_valid),
		.io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
		.io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
		.io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
		.io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
		.io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
		.io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data;
	assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid;
	assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode;
	assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param;
	assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size;
	assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source;
	assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address;
	assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask;
	assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data;
	assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready;
	assign bundleOut_0_a_q_clock = clock;
	assign bundleOut_0_a_q_reset = reset;
	assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid;
	assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param;
	assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size;
	assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source;
	assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address;
	assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask;
	assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data;
	assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready;
	assign bundleIn_0_d_q_clock = clock;
	assign bundleIn_0_d_q_reset = reset;
	assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid;
	assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign bundleIn_0_d_q_io_enq_bits_param = 2'h0;
	assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size;
	assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source;
	assign bundleIn_0_d_q_io_enq_bits_sink = 1'h0;
	assign bundleIn_0_d_q_io_enq_bits_denied = 1'h0;
	assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data;
	assign bundleIn_0_d_q_io_enq_bits_corrupt = 1'h0;
	assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready;
endmodule
module NonSyncResetSynchronizerPrimitiveShiftReg_d3 (
	clock,
	io_d,
	io_q
);
	input clock;
	input io_d;
	output wire io_q;
	reg sync_0;
	reg sync_1;
	reg sync_2;
	assign io_q = sync_0;
	always @(posedge clock) begin
		sync_0 <= sync_1;
		sync_1 <= sync_2;
		sync_2 <= io_d;
	end
endmodule
module SynchronizerShiftReg_w1_d3 (
	clock,
	io_d,
	io_q
);
	input clock;
	input io_d;
	output wire io_q;
	wire output_chain_clock;
	wire output_chain_io_d;
	wire output_chain_io_q;
	NonSyncResetSynchronizerPrimitiveShiftReg_d3 output_chain(
		.clock(output_chain_clock),
		.io_d(output_chain_io_d),
		.io_q(output_chain_io_q)
	);
	assign io_q = output_chain_io_q;
	assign output_chain_clock = clock;
	assign output_chain_io_d = io_d;
endmodule
module IntSyncAsyncCrossingSink (
	clock,
	auto_in_sync_0,
	auto_out_0
);
	input clock;
	input auto_in_sync_0;
	output wire auto_out_0;
	wire chain_clock;
	wire chain_io_d;
	wire chain_io_q;
	SynchronizerShiftReg_w1_d3 chain(
		.clock(chain_clock),
		.io_d(chain_io_d),
		.io_q(chain_io_q)
	);
	assign auto_out_0 = chain_io_q;
	assign chain_clock = clock;
	assign chain_io_d = auto_in_sync_0;
endmodule
module IntSyncSyncCrossingSink (
	auto_in_sync_0,
	auto_in_sync_1,
	auto_out_0,
	auto_out_1
);
	input auto_in_sync_0;
	input auto_in_sync_1;
	output wire auto_out_0;
	output wire auto_out_1;
	assign auto_out_0 = auto_in_sync_0;
	assign auto_out_1 = auto_in_sync_1;
endmodule
module IntSyncSyncCrossingSink_1 (
	auto_in_sync_0,
	auto_out_0
);
	input auto_in_sync_0;
	output wire auto_out_0;
	assign auto_out_0 = auto_in_sync_0;
endmodule
module AsyncResetRegVec_w1_i0 (
	clock,
	reset,
	io_d,
	io_q
);
	input clock;
	input reset;
	input io_d;
	output wire io_q;
	reg reg_;
	assign io_q = reg_;
	always @(posedge clock or posedge reset)
		if (reset)
			reg_ <= 1'h0;
		else
			reg_ <= io_d;
endmodule
module IntSyncCrossingSource_1 (
	clock,
	reset,
	auto_in_0,
	auto_out_sync_0
);
	input clock;
	input reset;
	input auto_in_0;
	output wire auto_out_sync_0;
	wire reg__clock;
	wire reg__reset;
	wire reg__io_d;
	wire reg__io_q;
	AsyncResetRegVec_w1_i0 reg_(
		.clock(reg__clock),
		.reset(reg__reset),
		.io_d(reg__io_d),
		.io_q(reg__io_q)
	);
	assign auto_out_sync_0 = reg__io_q;
	assign reg__clock = clock;
	assign reg__reset = reset;
	assign reg__io_d = auto_in_0;
endmodule
module TilePRCIDomain (
	auto_intsink_in_sync_0,
	auto_tile_reset_domain_tile_hartid_in,
	auto_int_out_clock_xing_out_2_sync_0,
	auto_int_out_clock_xing_out_1_sync_0,
	auto_int_out_clock_xing_out_0_sync_0,
	auto_int_in_clock_xing_in_1_sync_0,
	auto_int_in_clock_xing_in_0_sync_0,
	auto_int_in_clock_xing_in_0_sync_1,
	auto_tl_slave_clock_xing_in_a_ready,
	auto_tl_slave_clock_xing_in_a_valid,
	auto_tl_slave_clock_xing_in_a_bits_opcode,
	auto_tl_slave_clock_xing_in_a_bits_param,
	auto_tl_slave_clock_xing_in_a_bits_size,
	auto_tl_slave_clock_xing_in_a_bits_source,
	auto_tl_slave_clock_xing_in_a_bits_address,
	auto_tl_slave_clock_xing_in_a_bits_mask,
	auto_tl_slave_clock_xing_in_a_bits_data,
	auto_tl_slave_clock_xing_in_d_ready,
	auto_tl_slave_clock_xing_in_d_valid,
	auto_tl_slave_clock_xing_in_d_bits_opcode,
	auto_tl_slave_clock_xing_in_d_bits_param,
	auto_tl_slave_clock_xing_in_d_bits_size,
	auto_tl_slave_clock_xing_in_d_bits_source,
	auto_tl_slave_clock_xing_in_d_bits_sink,
	auto_tl_slave_clock_xing_in_d_bits_denied,
	auto_tl_slave_clock_xing_in_d_bits_data,
	auto_tl_slave_clock_xing_in_d_bits_corrupt,
	auto_tl_master_clock_xing_out_a_ready,
	auto_tl_master_clock_xing_out_a_valid,
	auto_tl_master_clock_xing_out_a_bits_opcode,
	auto_tl_master_clock_xing_out_a_bits_param,
	auto_tl_master_clock_xing_out_a_bits_size,
	auto_tl_master_clock_xing_out_a_bits_source,
	auto_tl_master_clock_xing_out_a_bits_address,
	auto_tl_master_clock_xing_out_a_bits_mask,
	auto_tl_master_clock_xing_out_a_bits_data,
	auto_tl_master_clock_xing_out_a_bits_corrupt,
	auto_tl_master_clock_xing_out_d_ready,
	auto_tl_master_clock_xing_out_d_valid,
	auto_tl_master_clock_xing_out_d_bits_opcode,
	auto_tl_master_clock_xing_out_d_bits_param,
	auto_tl_master_clock_xing_out_d_bits_size,
	auto_tl_master_clock_xing_out_d_bits_source,
	auto_tl_master_clock_xing_out_d_bits_sink,
	auto_tl_master_clock_xing_out_d_bits_denied,
	auto_tl_master_clock_xing_out_d_bits_data,
	auto_tl_master_clock_xing_out_d_bits_corrupt,
	auto_tap_clock_in_clock,
	auto_tap_clock_in_reset
);
	input auto_intsink_in_sync_0;
	input auto_tile_reset_domain_tile_hartid_in;
	output wire auto_int_out_clock_xing_out_2_sync_0;
	output wire auto_int_out_clock_xing_out_1_sync_0;
	output wire auto_int_out_clock_xing_out_0_sync_0;
	input auto_int_in_clock_xing_in_1_sync_0;
	input auto_int_in_clock_xing_in_0_sync_0;
	input auto_int_in_clock_xing_in_0_sync_1;
	output wire auto_tl_slave_clock_xing_in_a_ready;
	input auto_tl_slave_clock_xing_in_a_valid;
	input [2:0] auto_tl_slave_clock_xing_in_a_bits_opcode;
	input [2:0] auto_tl_slave_clock_xing_in_a_bits_param;
	input [2:0] auto_tl_slave_clock_xing_in_a_bits_size;
	input [2:0] auto_tl_slave_clock_xing_in_a_bits_source;
	input [31:0] auto_tl_slave_clock_xing_in_a_bits_address;
	input [3:0] auto_tl_slave_clock_xing_in_a_bits_mask;
	input [31:0] auto_tl_slave_clock_xing_in_a_bits_data;
	input auto_tl_slave_clock_xing_in_d_ready;
	output wire auto_tl_slave_clock_xing_in_d_valid;
	output wire [2:0] auto_tl_slave_clock_xing_in_d_bits_opcode;
	output wire [1:0] auto_tl_slave_clock_xing_in_d_bits_param;
	output wire [2:0] auto_tl_slave_clock_xing_in_d_bits_size;
	output wire [2:0] auto_tl_slave_clock_xing_in_d_bits_source;
	output wire auto_tl_slave_clock_xing_in_d_bits_sink;
	output wire auto_tl_slave_clock_xing_in_d_bits_denied;
	output wire [31:0] auto_tl_slave_clock_xing_in_d_bits_data;
	output wire auto_tl_slave_clock_xing_in_d_bits_corrupt;
	input auto_tl_master_clock_xing_out_a_ready;
	output wire auto_tl_master_clock_xing_out_a_valid;
	output wire [2:0] auto_tl_master_clock_xing_out_a_bits_opcode;
	output wire [2:0] auto_tl_master_clock_xing_out_a_bits_param;
	output wire [3:0] auto_tl_master_clock_xing_out_a_bits_size;
	output wire auto_tl_master_clock_xing_out_a_bits_source;
	output wire [31:0] auto_tl_master_clock_xing_out_a_bits_address;
	output wire [3:0] auto_tl_master_clock_xing_out_a_bits_mask;
	output wire [31:0] auto_tl_master_clock_xing_out_a_bits_data;
	output wire auto_tl_master_clock_xing_out_a_bits_corrupt;
	output wire auto_tl_master_clock_xing_out_d_ready;
	input auto_tl_master_clock_xing_out_d_valid;
	input [2:0] auto_tl_master_clock_xing_out_d_bits_opcode;
	input [1:0] auto_tl_master_clock_xing_out_d_bits_param;
	input [3:0] auto_tl_master_clock_xing_out_d_bits_size;
	input auto_tl_master_clock_xing_out_d_bits_source;
	input auto_tl_master_clock_xing_out_d_bits_sink;
	input auto_tl_master_clock_xing_out_d_bits_denied;
	input [31:0] auto_tl_master_clock_xing_out_d_bits_data;
	input auto_tl_master_clock_xing_out_d_bits_corrupt;
	input auto_tap_clock_in_clock;
	input auto_tap_clock_in_reset;
	wire tile_reset_domain_auto_tile_slave_in_a_ready;
	wire tile_reset_domain_auto_tile_slave_in_a_valid;
	wire [2:0] tile_reset_domain_auto_tile_slave_in_a_bits_opcode;
	wire [2:0] tile_reset_domain_auto_tile_slave_in_a_bits_param;
	wire [2:0] tile_reset_domain_auto_tile_slave_in_a_bits_size;
	wire [2:0] tile_reset_domain_auto_tile_slave_in_a_bits_source;
	wire [31:0] tile_reset_domain_auto_tile_slave_in_a_bits_address;
	wire [3:0] tile_reset_domain_auto_tile_slave_in_a_bits_mask;
	wire [31:0] tile_reset_domain_auto_tile_slave_in_a_bits_data;
	wire tile_reset_domain_auto_tile_slave_in_d_ready;
	wire tile_reset_domain_auto_tile_slave_in_d_valid;
	wire [2:0] tile_reset_domain_auto_tile_slave_in_d_bits_opcode;
	wire [2:0] tile_reset_domain_auto_tile_slave_in_d_bits_size;
	wire [2:0] tile_reset_domain_auto_tile_slave_in_d_bits_source;
	wire [31:0] tile_reset_domain_auto_tile_slave_in_d_bits_data;
	wire tile_reset_domain_auto_tile_wfi_out_0;
	wire tile_reset_domain_auto_tile_int_local_in_2_0;
	wire tile_reset_domain_auto_tile_int_local_in_1_0;
	wire tile_reset_domain_auto_tile_int_local_in_1_1;
	wire tile_reset_domain_auto_tile_int_local_in_0_0;
	wire tile_reset_domain_auto_tile_hartid_in;
	wire tile_reset_domain_auto_tile_tl_other_masters_out_a_ready;
	wire tile_reset_domain_auto_tile_tl_other_masters_out_a_valid;
	wire [2:0] tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_opcode;
	wire [2:0] tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_param;
	wire [3:0] tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_size;
	wire tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_source;
	wire [31:0] tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_address;
	wire [3:0] tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_mask;
	wire [31:0] tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_data;
	wire tile_reset_domain_auto_tile_tl_other_masters_out_d_ready;
	wire tile_reset_domain_auto_tile_tl_other_masters_out_d_valid;
	wire [2:0] tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_opcode;
	wire [1:0] tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_param;
	wire [3:0] tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_size;
	wire tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_source;
	wire tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_sink;
	wire tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_denied;
	wire [31:0] tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_data;
	wire tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_corrupt;
	wire tile_reset_domain_auto_clock_in_clock;
	wire tile_reset_domain_auto_clock_in_reset;
	wire clockNode_auto_in_clock;
	wire clockNode_auto_in_reset;
	wire clockNode_auto_out_clock;
	wire clockNode_auto_out_reset;
	wire buffer_auto_in_a_ready;
	wire buffer_auto_in_a_valid;
	wire [2:0] buffer_auto_in_a_bits_opcode;
	wire [2:0] buffer_auto_in_a_bits_param;
	wire [3:0] buffer_auto_in_a_bits_size;
	wire buffer_auto_in_a_bits_source;
	wire [31:0] buffer_auto_in_a_bits_address;
	wire [3:0] buffer_auto_in_a_bits_mask;
	wire [31:0] buffer_auto_in_a_bits_data;
	wire buffer_auto_in_d_ready;
	wire buffer_auto_in_d_valid;
	wire [2:0] buffer_auto_in_d_bits_opcode;
	wire [1:0] buffer_auto_in_d_bits_param;
	wire [3:0] buffer_auto_in_d_bits_size;
	wire buffer_auto_in_d_bits_source;
	wire buffer_auto_in_d_bits_sink;
	wire buffer_auto_in_d_bits_denied;
	wire [31:0] buffer_auto_in_d_bits_data;
	wire buffer_auto_in_d_bits_corrupt;
	wire buffer_auto_out_a_ready;
	wire buffer_auto_out_a_valid;
	wire [2:0] buffer_auto_out_a_bits_opcode;
	wire [2:0] buffer_auto_out_a_bits_param;
	wire [3:0] buffer_auto_out_a_bits_size;
	wire buffer_auto_out_a_bits_source;
	wire [31:0] buffer_auto_out_a_bits_address;
	wire [3:0] buffer_auto_out_a_bits_mask;
	wire [31:0] buffer_auto_out_a_bits_data;
	wire buffer_auto_out_d_ready;
	wire buffer_auto_out_d_valid;
	wire [2:0] buffer_auto_out_d_bits_opcode;
	wire [1:0] buffer_auto_out_d_bits_param;
	wire [3:0] buffer_auto_out_d_bits_size;
	wire buffer_auto_out_d_bits_source;
	wire buffer_auto_out_d_bits_sink;
	wire buffer_auto_out_d_bits_denied;
	wire [31:0] buffer_auto_out_d_bits_data;
	wire buffer_auto_out_d_bits_corrupt;
	wire buffer_1_clock;
	wire buffer_1_reset;
	wire buffer_1_auto_in_a_ready;
	wire buffer_1_auto_in_a_valid;
	wire [2:0] buffer_1_auto_in_a_bits_opcode;
	wire [2:0] buffer_1_auto_in_a_bits_param;
	wire [3:0] buffer_1_auto_in_a_bits_size;
	wire buffer_1_auto_in_a_bits_source;
	wire [31:0] buffer_1_auto_in_a_bits_address;
	wire [3:0] buffer_1_auto_in_a_bits_mask;
	wire [31:0] buffer_1_auto_in_a_bits_data;
	wire buffer_1_auto_in_d_ready;
	wire buffer_1_auto_in_d_valid;
	wire [2:0] buffer_1_auto_in_d_bits_opcode;
	wire [1:0] buffer_1_auto_in_d_bits_param;
	wire [3:0] buffer_1_auto_in_d_bits_size;
	wire buffer_1_auto_in_d_bits_source;
	wire buffer_1_auto_in_d_bits_sink;
	wire buffer_1_auto_in_d_bits_denied;
	wire [31:0] buffer_1_auto_in_d_bits_data;
	wire buffer_1_auto_in_d_bits_corrupt;
	wire buffer_1_auto_out_a_ready;
	wire buffer_1_auto_out_a_valid;
	wire [2:0] buffer_1_auto_out_a_bits_opcode;
	wire [2:0] buffer_1_auto_out_a_bits_param;
	wire [3:0] buffer_1_auto_out_a_bits_size;
	wire buffer_1_auto_out_a_bits_source;
	wire [31:0] buffer_1_auto_out_a_bits_address;
	wire [3:0] buffer_1_auto_out_a_bits_mask;
	wire [31:0] buffer_1_auto_out_a_bits_data;
	wire buffer_1_auto_out_a_bits_corrupt;
	wire buffer_1_auto_out_d_ready;
	wire buffer_1_auto_out_d_valid;
	wire [2:0] buffer_1_auto_out_d_bits_opcode;
	wire [1:0] buffer_1_auto_out_d_bits_param;
	wire [3:0] buffer_1_auto_out_d_bits_size;
	wire buffer_1_auto_out_d_bits_source;
	wire buffer_1_auto_out_d_bits_sink;
	wire buffer_1_auto_out_d_bits_denied;
	wire [31:0] buffer_1_auto_out_d_bits_data;
	wire buffer_1_auto_out_d_bits_corrupt;
	wire buffer_2_auto_in_a_ready;
	wire buffer_2_auto_in_a_valid;
	wire [2:0] buffer_2_auto_in_a_bits_opcode;
	wire [2:0] buffer_2_auto_in_a_bits_param;
	wire [2:0] buffer_2_auto_in_a_bits_size;
	wire [2:0] buffer_2_auto_in_a_bits_source;
	wire [31:0] buffer_2_auto_in_a_bits_address;
	wire [3:0] buffer_2_auto_in_a_bits_mask;
	wire [31:0] buffer_2_auto_in_a_bits_data;
	wire buffer_2_auto_in_d_ready;
	wire buffer_2_auto_in_d_valid;
	wire [2:0] buffer_2_auto_in_d_bits_opcode;
	wire [2:0] buffer_2_auto_in_d_bits_size;
	wire [2:0] buffer_2_auto_in_d_bits_source;
	wire [31:0] buffer_2_auto_in_d_bits_data;
	wire buffer_2_auto_out_a_ready;
	wire buffer_2_auto_out_a_valid;
	wire [2:0] buffer_2_auto_out_a_bits_opcode;
	wire [2:0] buffer_2_auto_out_a_bits_param;
	wire [2:0] buffer_2_auto_out_a_bits_size;
	wire [2:0] buffer_2_auto_out_a_bits_source;
	wire [31:0] buffer_2_auto_out_a_bits_address;
	wire [3:0] buffer_2_auto_out_a_bits_mask;
	wire [31:0] buffer_2_auto_out_a_bits_data;
	wire buffer_2_auto_out_d_ready;
	wire buffer_2_auto_out_d_valid;
	wire [2:0] buffer_2_auto_out_d_bits_opcode;
	wire [2:0] buffer_2_auto_out_d_bits_size;
	wire [2:0] buffer_2_auto_out_d_bits_source;
	wire [31:0] buffer_2_auto_out_d_bits_data;
	wire buffer_3_clock;
	wire buffer_3_reset;
	wire buffer_3_auto_in_a_ready;
	wire buffer_3_auto_in_a_valid;
	wire [2:0] buffer_3_auto_in_a_bits_opcode;
	wire [2:0] buffer_3_auto_in_a_bits_param;
	wire [2:0] buffer_3_auto_in_a_bits_size;
	wire [2:0] buffer_3_auto_in_a_bits_source;
	wire [31:0] buffer_3_auto_in_a_bits_address;
	wire [3:0] buffer_3_auto_in_a_bits_mask;
	wire [31:0] buffer_3_auto_in_a_bits_data;
	wire buffer_3_auto_in_d_ready;
	wire buffer_3_auto_in_d_valid;
	wire [2:0] buffer_3_auto_in_d_bits_opcode;
	wire [1:0] buffer_3_auto_in_d_bits_param;
	wire [2:0] buffer_3_auto_in_d_bits_size;
	wire [2:0] buffer_3_auto_in_d_bits_source;
	wire buffer_3_auto_in_d_bits_sink;
	wire buffer_3_auto_in_d_bits_denied;
	wire [31:0] buffer_3_auto_in_d_bits_data;
	wire buffer_3_auto_in_d_bits_corrupt;
	wire buffer_3_auto_out_a_ready;
	wire buffer_3_auto_out_a_valid;
	wire [2:0] buffer_3_auto_out_a_bits_opcode;
	wire [2:0] buffer_3_auto_out_a_bits_param;
	wire [2:0] buffer_3_auto_out_a_bits_size;
	wire [2:0] buffer_3_auto_out_a_bits_source;
	wire [31:0] buffer_3_auto_out_a_bits_address;
	wire [3:0] buffer_3_auto_out_a_bits_mask;
	wire [31:0] buffer_3_auto_out_a_bits_data;
	wire buffer_3_auto_out_d_ready;
	wire buffer_3_auto_out_d_valid;
	wire [2:0] buffer_3_auto_out_d_bits_opcode;
	wire [2:0] buffer_3_auto_out_d_bits_size;
	wire [2:0] buffer_3_auto_out_d_bits_source;
	wire [31:0] buffer_3_auto_out_d_bits_data;
	wire intsink_clock;
	wire intsink_auto_in_sync_0;
	wire intsink_auto_out_0;
	wire intsink_1_auto_in_sync_0;
	wire intsink_1_auto_in_sync_1;
	wire intsink_1_auto_out_0;
	wire intsink_1_auto_out_1;
	wire intsink_2_auto_in_sync_0;
	wire intsink_2_auto_out_0;
	wire intsource_1_clock;
	wire intsource_1_reset;
	wire intsource_1_auto_in_0;
	wire intsource_1_auto_out_sync_0;
	wire intsource_2_clock;
	wire intsource_2_reset;
	wire intsource_2_auto_in_0;
	wire intsource_2_auto_out_sync_0;
	wire intsource_3_clock;
	wire intsource_3_reset;
	wire intsource_3_auto_in_0;
	wire intsource_3_auto_out_sync_0;
	TileResetDomain tile_reset_domain(
		.auto_tile_slave_in_a_ready(tile_reset_domain_auto_tile_slave_in_a_ready),
		.auto_tile_slave_in_a_valid(tile_reset_domain_auto_tile_slave_in_a_valid),
		.auto_tile_slave_in_a_bits_opcode(tile_reset_domain_auto_tile_slave_in_a_bits_opcode),
		.auto_tile_slave_in_a_bits_param(tile_reset_domain_auto_tile_slave_in_a_bits_param),
		.auto_tile_slave_in_a_bits_size(tile_reset_domain_auto_tile_slave_in_a_bits_size),
		.auto_tile_slave_in_a_bits_source(tile_reset_domain_auto_tile_slave_in_a_bits_source),
		.auto_tile_slave_in_a_bits_address(tile_reset_domain_auto_tile_slave_in_a_bits_address),
		.auto_tile_slave_in_a_bits_mask(tile_reset_domain_auto_tile_slave_in_a_bits_mask),
		.auto_tile_slave_in_a_bits_data(tile_reset_domain_auto_tile_slave_in_a_bits_data),
		.auto_tile_slave_in_d_ready(tile_reset_domain_auto_tile_slave_in_d_ready),
		.auto_tile_slave_in_d_valid(tile_reset_domain_auto_tile_slave_in_d_valid),
		.auto_tile_slave_in_d_bits_opcode(tile_reset_domain_auto_tile_slave_in_d_bits_opcode),
		.auto_tile_slave_in_d_bits_size(tile_reset_domain_auto_tile_slave_in_d_bits_size),
		.auto_tile_slave_in_d_bits_source(tile_reset_domain_auto_tile_slave_in_d_bits_source),
		.auto_tile_slave_in_d_bits_data(tile_reset_domain_auto_tile_slave_in_d_bits_data),
		.auto_tile_wfi_out_0(tile_reset_domain_auto_tile_wfi_out_0),
		.auto_tile_int_local_in_2_0(tile_reset_domain_auto_tile_int_local_in_2_0),
		.auto_tile_int_local_in_1_0(tile_reset_domain_auto_tile_int_local_in_1_0),
		.auto_tile_int_local_in_1_1(tile_reset_domain_auto_tile_int_local_in_1_1),
		.auto_tile_int_local_in_0_0(tile_reset_domain_auto_tile_int_local_in_0_0),
		.auto_tile_hartid_in(tile_reset_domain_auto_tile_hartid_in),
		.auto_tile_tl_other_masters_out_a_ready(tile_reset_domain_auto_tile_tl_other_masters_out_a_ready),
		.auto_tile_tl_other_masters_out_a_valid(tile_reset_domain_auto_tile_tl_other_masters_out_a_valid),
		.auto_tile_tl_other_masters_out_a_bits_opcode(tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_opcode),
		.auto_tile_tl_other_masters_out_a_bits_param(tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_param),
		.auto_tile_tl_other_masters_out_a_bits_size(tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_size),
		.auto_tile_tl_other_masters_out_a_bits_source(tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_source),
		.auto_tile_tl_other_masters_out_a_bits_address(tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_address),
		.auto_tile_tl_other_masters_out_a_bits_mask(tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_mask),
		.auto_tile_tl_other_masters_out_a_bits_data(tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_data),
		.auto_tile_tl_other_masters_out_d_ready(tile_reset_domain_auto_tile_tl_other_masters_out_d_ready),
		.auto_tile_tl_other_masters_out_d_valid(tile_reset_domain_auto_tile_tl_other_masters_out_d_valid),
		.auto_tile_tl_other_masters_out_d_bits_opcode(tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_opcode),
		.auto_tile_tl_other_masters_out_d_bits_param(tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_param),
		.auto_tile_tl_other_masters_out_d_bits_size(tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_size),
		.auto_tile_tl_other_masters_out_d_bits_source(tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_source),
		.auto_tile_tl_other_masters_out_d_bits_sink(tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_sink),
		.auto_tile_tl_other_masters_out_d_bits_denied(tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_denied),
		.auto_tile_tl_other_masters_out_d_bits_data(tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_data),
		.auto_tile_tl_other_masters_out_d_bits_corrupt(tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_corrupt),
		.auto_clock_in_clock(tile_reset_domain_auto_clock_in_clock),
		.auto_clock_in_reset(tile_reset_domain_auto_clock_in_reset)
	);
	FixedClockBroadcast_4 clockNode(
		.auto_in_clock(clockNode_auto_in_clock),
		.auto_in_reset(clockNode_auto_in_reset),
		.auto_out_clock(clockNode_auto_out_clock),
		.auto_out_reset(clockNode_auto_out_reset)
	);
	TLBuffer_13 buffer(
		.auto_in_a_ready(buffer_auto_in_a_ready),
		.auto_in_a_valid(buffer_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_auto_in_a_bits_data),
		.auto_in_d_ready(buffer_auto_in_d_ready),
		.auto_in_d_valid(buffer_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_auto_out_a_ready),
		.auto_out_a_valid(buffer_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_auto_out_a_bits_data),
		.auto_out_d_ready(buffer_auto_out_d_ready),
		.auto_out_d_valid(buffer_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(buffer_auto_out_d_bits_param),
		.auto_out_d_bits_size(buffer_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_auto_out_d_bits_source),
		.auto_out_d_bits_sink(buffer_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
		.auto_out_d_bits_data(buffer_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt)
	);
	TLBuffer_14 buffer_1(
		.clock(buffer_1_clock),
		.reset(buffer_1_reset),
		.auto_in_a_ready(buffer_1_auto_in_a_ready),
		.auto_in_a_valid(buffer_1_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_1_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_1_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_1_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_1_auto_in_a_bits_data),
		.auto_in_d_ready(buffer_1_auto_in_d_ready),
		.auto_in_d_valid(buffer_1_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_1_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_1_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_1_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_1_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_1_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_1_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_1_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_1_auto_out_a_ready),
		.auto_out_a_valid(buffer_1_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_1_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_1_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_1_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_1_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_1_auto_out_d_ready),
		.auto_out_d_valid(buffer_1_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(buffer_1_auto_out_d_bits_param),
		.auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
		.auto_out_d_bits_sink(buffer_1_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
		.auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt)
	);
	TLBuffer_15 buffer_2(
		.auto_in_a_ready(buffer_2_auto_in_a_ready),
		.auto_in_a_valid(buffer_2_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_2_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_2_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_2_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_2_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_2_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_2_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_2_auto_in_a_bits_data),
		.auto_in_d_ready(buffer_2_auto_in_d_ready),
		.auto_in_d_valid(buffer_2_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_2_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(buffer_2_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_2_auto_in_d_bits_source),
		.auto_in_d_bits_data(buffer_2_auto_in_d_bits_data),
		.auto_out_a_ready(buffer_2_auto_out_a_ready),
		.auto_out_a_valid(buffer_2_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_2_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_2_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_2_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_2_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_2_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_2_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_2_auto_out_a_bits_data),
		.auto_out_d_ready(buffer_2_auto_out_d_ready),
		.auto_out_d_valid(buffer_2_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_2_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(buffer_2_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_2_auto_out_d_bits_source),
		.auto_out_d_bits_data(buffer_2_auto_out_d_bits_data)
	);
	TLBuffer_16 buffer_3(
		.clock(buffer_3_clock),
		.reset(buffer_3_reset),
		.auto_in_a_ready(buffer_3_auto_in_a_ready),
		.auto_in_a_valid(buffer_3_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_3_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_3_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_3_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_3_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_3_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_3_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_3_auto_in_a_bits_data),
		.auto_in_d_ready(buffer_3_auto_in_d_ready),
		.auto_in_d_valid(buffer_3_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_3_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_3_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_3_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_3_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_3_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_3_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_3_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_3_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_3_auto_out_a_ready),
		.auto_out_a_valid(buffer_3_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_3_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_3_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_3_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_3_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_3_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_3_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_3_auto_out_a_bits_data),
		.auto_out_d_ready(buffer_3_auto_out_d_ready),
		.auto_out_d_valid(buffer_3_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_3_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(buffer_3_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_3_auto_out_d_bits_source),
		.auto_out_d_bits_data(buffer_3_auto_out_d_bits_data)
	);
	IntSyncAsyncCrossingSink intsink(
		.clock(intsink_clock),
		.auto_in_sync_0(intsink_auto_in_sync_0),
		.auto_out_0(intsink_auto_out_0)
	);
	IntSyncSyncCrossingSink intsink_1(
		.auto_in_sync_0(intsink_1_auto_in_sync_0),
		.auto_in_sync_1(intsink_1_auto_in_sync_1),
		.auto_out_0(intsink_1_auto_out_0),
		.auto_out_1(intsink_1_auto_out_1)
	);
	IntSyncSyncCrossingSink_1 intsink_2(
		.auto_in_sync_0(intsink_2_auto_in_sync_0),
		.auto_out_0(intsink_2_auto_out_0)
	);
	IntSyncCrossingSource_1 intsource_1(
		.clock(intsource_1_clock),
		.reset(intsource_1_reset),
		.auto_in_0(intsource_1_auto_in_0),
		.auto_out_sync_0(intsource_1_auto_out_sync_0)
	);
	IntSyncCrossingSource_1 intsource_2(
		.clock(intsource_2_clock),
		.reset(intsource_2_reset),
		.auto_in_0(intsource_2_auto_in_0),
		.auto_out_sync_0(intsource_2_auto_out_sync_0)
	);
	IntSyncCrossingSource_1 intsource_3(
		.clock(intsource_3_clock),
		.reset(intsource_3_reset),
		.auto_in_0(intsource_3_auto_in_0),
		.auto_out_sync_0(intsource_3_auto_out_sync_0)
	);
	assign auto_int_out_clock_xing_out_2_sync_0 = intsource_3_auto_out_sync_0;
	assign auto_int_out_clock_xing_out_1_sync_0 = intsource_2_auto_out_sync_0;
	assign auto_int_out_clock_xing_out_0_sync_0 = intsource_1_auto_out_sync_0;
	assign auto_tl_slave_clock_xing_in_a_ready = buffer_3_auto_in_a_ready;
	assign auto_tl_slave_clock_xing_in_d_valid = buffer_3_auto_in_d_valid;
	assign auto_tl_slave_clock_xing_in_d_bits_opcode = buffer_3_auto_in_d_bits_opcode;
	assign auto_tl_slave_clock_xing_in_d_bits_param = buffer_3_auto_in_d_bits_param;
	assign auto_tl_slave_clock_xing_in_d_bits_size = buffer_3_auto_in_d_bits_size;
	assign auto_tl_slave_clock_xing_in_d_bits_source = buffer_3_auto_in_d_bits_source;
	assign auto_tl_slave_clock_xing_in_d_bits_sink = buffer_3_auto_in_d_bits_sink;
	assign auto_tl_slave_clock_xing_in_d_bits_denied = buffer_3_auto_in_d_bits_denied;
	assign auto_tl_slave_clock_xing_in_d_bits_data = buffer_3_auto_in_d_bits_data;
	assign auto_tl_slave_clock_xing_in_d_bits_corrupt = buffer_3_auto_in_d_bits_corrupt;
	assign auto_tl_master_clock_xing_out_a_valid = buffer_1_auto_out_a_valid;
	assign auto_tl_master_clock_xing_out_a_bits_opcode = buffer_1_auto_out_a_bits_opcode;
	assign auto_tl_master_clock_xing_out_a_bits_param = buffer_1_auto_out_a_bits_param;
	assign auto_tl_master_clock_xing_out_a_bits_size = buffer_1_auto_out_a_bits_size;
	assign auto_tl_master_clock_xing_out_a_bits_source = buffer_1_auto_out_a_bits_source;
	assign auto_tl_master_clock_xing_out_a_bits_address = buffer_1_auto_out_a_bits_address;
	assign auto_tl_master_clock_xing_out_a_bits_mask = buffer_1_auto_out_a_bits_mask;
	assign auto_tl_master_clock_xing_out_a_bits_data = buffer_1_auto_out_a_bits_data;
	assign auto_tl_master_clock_xing_out_a_bits_corrupt = buffer_1_auto_out_a_bits_corrupt;
	assign auto_tl_master_clock_xing_out_d_ready = buffer_1_auto_out_d_ready;
	assign tile_reset_domain_auto_tile_slave_in_a_valid = buffer_2_auto_out_a_valid;
	assign tile_reset_domain_auto_tile_slave_in_a_bits_opcode = buffer_2_auto_out_a_bits_opcode;
	assign tile_reset_domain_auto_tile_slave_in_a_bits_param = buffer_2_auto_out_a_bits_param;
	assign tile_reset_domain_auto_tile_slave_in_a_bits_size = buffer_2_auto_out_a_bits_size;
	assign tile_reset_domain_auto_tile_slave_in_a_bits_source = buffer_2_auto_out_a_bits_source;
	assign tile_reset_domain_auto_tile_slave_in_a_bits_address = buffer_2_auto_out_a_bits_address;
	assign tile_reset_domain_auto_tile_slave_in_a_bits_mask = buffer_2_auto_out_a_bits_mask;
	assign tile_reset_domain_auto_tile_slave_in_a_bits_data = buffer_2_auto_out_a_bits_data;
	assign tile_reset_domain_auto_tile_slave_in_d_ready = buffer_2_auto_out_d_ready;
	assign tile_reset_domain_auto_tile_int_local_in_2_0 = intsink_2_auto_out_0;
	assign tile_reset_domain_auto_tile_int_local_in_1_0 = intsink_1_auto_out_0;
	assign tile_reset_domain_auto_tile_int_local_in_1_1 = intsink_1_auto_out_1;
	assign tile_reset_domain_auto_tile_int_local_in_0_0 = intsink_auto_out_0;
	assign tile_reset_domain_auto_tile_hartid_in = auto_tile_reset_domain_tile_hartid_in;
	assign tile_reset_domain_auto_tile_tl_other_masters_out_a_ready = buffer_auto_in_a_ready;
	assign tile_reset_domain_auto_tile_tl_other_masters_out_d_valid = buffer_auto_in_d_valid;
	assign tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_opcode = buffer_auto_in_d_bits_opcode;
	assign tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_param = buffer_auto_in_d_bits_param;
	assign tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_size = buffer_auto_in_d_bits_size;
	assign tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_source = buffer_auto_in_d_bits_source;
	assign tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_sink = buffer_auto_in_d_bits_sink;
	assign tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_denied = buffer_auto_in_d_bits_denied;
	assign tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_data = buffer_auto_in_d_bits_data;
	assign tile_reset_domain_auto_tile_tl_other_masters_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt;
	assign tile_reset_domain_auto_clock_in_clock = clockNode_auto_out_clock;
	assign tile_reset_domain_auto_clock_in_reset = clockNode_auto_out_reset;
	assign clockNode_auto_in_clock = auto_tap_clock_in_clock;
	assign clockNode_auto_in_reset = auto_tap_clock_in_reset;
	assign buffer_auto_in_a_valid = tile_reset_domain_auto_tile_tl_other_masters_out_a_valid;
	assign buffer_auto_in_a_bits_opcode = tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_opcode;
	assign buffer_auto_in_a_bits_param = tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_param;
	assign buffer_auto_in_a_bits_size = tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_size;
	assign buffer_auto_in_a_bits_source = tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_source;
	assign buffer_auto_in_a_bits_address = tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_address;
	assign buffer_auto_in_a_bits_mask = tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_mask;
	assign buffer_auto_in_a_bits_data = tile_reset_domain_auto_tile_tl_other_masters_out_a_bits_data;
	assign buffer_auto_in_d_ready = tile_reset_domain_auto_tile_tl_other_masters_out_d_ready;
	assign buffer_auto_out_a_ready = buffer_1_auto_in_a_ready;
	assign buffer_auto_out_d_valid = buffer_1_auto_in_d_valid;
	assign buffer_auto_out_d_bits_opcode = buffer_1_auto_in_d_bits_opcode;
	assign buffer_auto_out_d_bits_param = buffer_1_auto_in_d_bits_param;
	assign buffer_auto_out_d_bits_size = buffer_1_auto_in_d_bits_size;
	assign buffer_auto_out_d_bits_source = buffer_1_auto_in_d_bits_source;
	assign buffer_auto_out_d_bits_sink = buffer_1_auto_in_d_bits_sink;
	assign buffer_auto_out_d_bits_denied = buffer_1_auto_in_d_bits_denied;
	assign buffer_auto_out_d_bits_data = buffer_1_auto_in_d_bits_data;
	assign buffer_auto_out_d_bits_corrupt = buffer_1_auto_in_d_bits_corrupt;
	assign buffer_1_clock = auto_tap_clock_in_clock;
	assign buffer_1_reset = auto_tap_clock_in_reset;
	assign buffer_1_auto_in_a_valid = buffer_auto_out_a_valid;
	assign buffer_1_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode;
	assign buffer_1_auto_in_a_bits_param = buffer_auto_out_a_bits_param;
	assign buffer_1_auto_in_a_bits_size = buffer_auto_out_a_bits_size;
	assign buffer_1_auto_in_a_bits_source = buffer_auto_out_a_bits_source;
	assign buffer_1_auto_in_a_bits_address = buffer_auto_out_a_bits_address;
	assign buffer_1_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask;
	assign buffer_1_auto_in_a_bits_data = buffer_auto_out_a_bits_data;
	assign buffer_1_auto_in_d_ready = buffer_auto_out_d_ready;
	assign buffer_1_auto_out_a_ready = auto_tl_master_clock_xing_out_a_ready;
	assign buffer_1_auto_out_d_valid = auto_tl_master_clock_xing_out_d_valid;
	assign buffer_1_auto_out_d_bits_opcode = auto_tl_master_clock_xing_out_d_bits_opcode;
	assign buffer_1_auto_out_d_bits_param = auto_tl_master_clock_xing_out_d_bits_param;
	assign buffer_1_auto_out_d_bits_size = auto_tl_master_clock_xing_out_d_bits_size;
	assign buffer_1_auto_out_d_bits_source = auto_tl_master_clock_xing_out_d_bits_source;
	assign buffer_1_auto_out_d_bits_sink = auto_tl_master_clock_xing_out_d_bits_sink;
	assign buffer_1_auto_out_d_bits_denied = auto_tl_master_clock_xing_out_d_bits_denied;
	assign buffer_1_auto_out_d_bits_data = auto_tl_master_clock_xing_out_d_bits_data;
	assign buffer_1_auto_out_d_bits_corrupt = auto_tl_master_clock_xing_out_d_bits_corrupt;
	assign buffer_2_auto_in_a_valid = buffer_3_auto_out_a_valid;
	assign buffer_2_auto_in_a_bits_opcode = buffer_3_auto_out_a_bits_opcode;
	assign buffer_2_auto_in_a_bits_param = buffer_3_auto_out_a_bits_param;
	assign buffer_2_auto_in_a_bits_size = buffer_3_auto_out_a_bits_size;
	assign buffer_2_auto_in_a_bits_source = buffer_3_auto_out_a_bits_source;
	assign buffer_2_auto_in_a_bits_address = buffer_3_auto_out_a_bits_address;
	assign buffer_2_auto_in_a_bits_mask = buffer_3_auto_out_a_bits_mask;
	assign buffer_2_auto_in_a_bits_data = buffer_3_auto_out_a_bits_data;
	assign buffer_2_auto_in_d_ready = buffer_3_auto_out_d_ready;
	assign buffer_2_auto_out_a_ready = tile_reset_domain_auto_tile_slave_in_a_ready;
	assign buffer_2_auto_out_d_valid = tile_reset_domain_auto_tile_slave_in_d_valid;
	assign buffer_2_auto_out_d_bits_opcode = tile_reset_domain_auto_tile_slave_in_d_bits_opcode;
	assign buffer_2_auto_out_d_bits_size = tile_reset_domain_auto_tile_slave_in_d_bits_size;
	assign buffer_2_auto_out_d_bits_source = tile_reset_domain_auto_tile_slave_in_d_bits_source;
	assign buffer_2_auto_out_d_bits_data = tile_reset_domain_auto_tile_slave_in_d_bits_data;
	assign buffer_3_clock = auto_tap_clock_in_clock;
	assign buffer_3_reset = auto_tap_clock_in_reset;
	assign buffer_3_auto_in_a_valid = auto_tl_slave_clock_xing_in_a_valid;
	assign buffer_3_auto_in_a_bits_opcode = auto_tl_slave_clock_xing_in_a_bits_opcode;
	assign buffer_3_auto_in_a_bits_param = auto_tl_slave_clock_xing_in_a_bits_param;
	assign buffer_3_auto_in_a_bits_size = auto_tl_slave_clock_xing_in_a_bits_size;
	assign buffer_3_auto_in_a_bits_source = auto_tl_slave_clock_xing_in_a_bits_source;
	assign buffer_3_auto_in_a_bits_address = auto_tl_slave_clock_xing_in_a_bits_address;
	assign buffer_3_auto_in_a_bits_mask = auto_tl_slave_clock_xing_in_a_bits_mask;
	assign buffer_3_auto_in_a_bits_data = auto_tl_slave_clock_xing_in_a_bits_data;
	assign buffer_3_auto_in_d_ready = auto_tl_slave_clock_xing_in_d_ready;
	assign buffer_3_auto_out_a_ready = buffer_2_auto_in_a_ready;
	assign buffer_3_auto_out_d_valid = buffer_2_auto_in_d_valid;
	assign buffer_3_auto_out_d_bits_opcode = buffer_2_auto_in_d_bits_opcode;
	assign buffer_3_auto_out_d_bits_size = buffer_2_auto_in_d_bits_size;
	assign buffer_3_auto_out_d_bits_source = buffer_2_auto_in_d_bits_source;
	assign buffer_3_auto_out_d_bits_data = buffer_2_auto_in_d_bits_data;
	assign intsink_clock = auto_tap_clock_in_clock;
	assign intsink_auto_in_sync_0 = auto_intsink_in_sync_0;
	assign intsink_1_auto_in_sync_0 = auto_int_in_clock_xing_in_0_sync_0;
	assign intsink_1_auto_in_sync_1 = auto_int_in_clock_xing_in_0_sync_1;
	assign intsink_2_auto_in_sync_0 = auto_int_in_clock_xing_in_1_sync_0;
	assign intsource_1_clock = auto_tap_clock_in_clock;
	assign intsource_1_reset = auto_tap_clock_in_reset;
	assign intsource_1_auto_in_0 = 1'h0;
	assign intsource_2_clock = auto_tap_clock_in_clock;
	assign intsource_2_reset = auto_tap_clock_in_reset;
	assign intsource_2_auto_in_0 = tile_reset_domain_auto_tile_wfi_out_0;
	assign intsource_3_clock = auto_tap_clock_in_clock;
	assign intsource_3_reset = auto_tap_clock_in_reset;
	assign intsource_3_auto_in_0 = 1'h0;
endmodule
module TLMonitor_34 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [1:0] io_in_a_bits_size;
	input [7:0] io_in_a_bits_source;
	input [27:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_size;
	input [7:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_4 = io_in_a_bits_source <= 8'h9f;
	wire [4:0] _is_aligned_mask_T_1 = 5'h03 << io_in_a_bits_size;
	wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0];
	wire [27:0] _GEN_71 = {26'd0, is_aligned_mask};
	wire [27:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 28'h0000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 2'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_10 = ~_source_ok_T_4;
	wire _T_20 = io_in_a_bits_opcode == 3'h6;
	wire [27:0] _T_33 = io_in_a_bits_address ^ 28'hc000000;
	wire [28:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [28:0] _T_36 = $signed(_T_34) & -29'sh04000000;
	wire _T_37 = $signed(_T_36) == 29'sh00000000;
	wire _T_69 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_73 = ~io_in_a_bits_mask;
	wire _T_74 = _T_73 == 4'h0;
	wire _T_78 = ~io_in_a_bits_corrupt;
	wire _T_82 = io_in_a_bits_opcode == 3'h7;
	wire _T_135 = io_in_a_bits_param != 3'h0;
	wire _T_148 = io_in_a_bits_opcode == 3'h4;
	wire _T_164 = io_in_a_bits_size <= 2'h2;
	wire _T_172 = _T_164 & _T_37;
	wire _T_183 = io_in_a_bits_param == 3'h0;
	wire _T_187 = io_in_a_bits_mask == mask;
	wire _T_195 = io_in_a_bits_opcode == 3'h0;
	wire _T_218 = _source_ok_T_4 & _T_172;
	wire _T_236 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_273 = ~mask;
	wire [3:0] _T_274 = io_in_a_bits_mask & _T_273;
	wire _T_275 = _T_274 == 4'h0;
	wire _T_279 = io_in_a_bits_opcode == 3'h2;
	wire _T_309 = io_in_a_bits_param <= 3'h4;
	wire _T_317 = io_in_a_bits_opcode == 3'h3;
	wire _T_347 = io_in_a_bits_param <= 3'h3;
	wire _T_355 = io_in_a_bits_opcode == 3'h5;
	wire _T_385 = io_in_a_bits_param <= 3'h1;
	wire _T_397 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_10 = io_in_d_bits_source <= 8'h9f;
	wire _T_401 = io_in_d_bits_opcode == 3'h6;
	wire _T_405 = io_in_d_bits_size >= 2'h2;
	wire _T_421 = io_in_d_bits_opcode == 3'h4;
	wire _T_449 = io_in_d_bits_opcode == 3'h5;
	wire _T_478 = io_in_d_bits_opcode == 3'h0;
	wire _T_495 = io_in_d_bits_opcode == 3'h1;
	wire _T_513 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [1:0] size;
	reg [7:0] source;
	reg [27:0] address;
	wire _T_543 = io_in_a_valid & ~a_first;
	wire _T_544 = io_in_a_bits_opcode == opcode;
	wire _T_548 = io_in_a_bits_param == param;
	wire _T_552 = io_in_a_bits_size == size;
	wire _T_556 = io_in_a_bits_source == source;
	wire _T_560 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] size_1;
	reg [7:0] source_1;
	wire _T_567 = io_in_d_valid & ~d_first;
	wire _T_568 = io_in_d_bits_opcode == opcode_1;
	wire _T_576 = io_in_d_bits_size == size_1;
	wire _T_580 = io_in_d_bits_source == source_1;
	reg [159:0] inflight;
	reg [639:0] inflight_opcodes;
	reg [639:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [10:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [639:0] _GEN_73 = {624'd0, _a_opcode_lookup_T_5};
	wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [639:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[639:1]};
	wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [639:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[639:1]};
	wire _T_594 = io_in_a_valid & a_first_1;
	wire [255:0] _a_set_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_a_bits_source;
	wire [255:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire _T_597 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1;
	wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [10:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [2050:0] _GEN_1 = {2047'd0, a_opcodes_set_interm};
	wire [2050:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? _a_sizes_set_interm_T_1 : 3'h0);
	wire [2049:0] _GEN_2 = {2047'd0, a_sizes_set_interm};
	wire [2049:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [159:0] _T_599 = inflight >> io_in_a_bits_source;
	wire _T_601 = ~_T_599[0];
	wire [255:0] _GEN_16 = (a_first_done & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2050:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 2051'h0);
	wire [2049:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 2050'h0);
	wire _T_605 = io_in_d_valid & d_first_1;
	wire _T_607 = ~_T_401;
	wire _T_608 = (io_in_d_valid & d_first_1) & ~_T_401;
	wire [255:0] _d_clr_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_d_bits_source;
	wire [255:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_401 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_3 = {2047'd0, _a_opcode_lookup_T_5};
	wire [2062:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [255:0] _GEN_22 = ((d_first_done & d_first_1) & _T_607 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_23 = ((d_first_done & d_first_1) & _T_607 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_594 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [159:0] _T_618 = inflight >> io_in_d_bits_source;
	wire _T_620 = _T_618[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_625 = io_in_d_bits_opcode == _GEN_40;
	wire _T_626 = (io_in_d_bits_opcode == _GEN_32) | _T_625;
	wire _T_630 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_637 = io_in_d_bits_opcode == _GEN_56;
	wire _T_638 = (io_in_d_bits_opcode == _GEN_48) | _T_637;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {2'd0, io_in_d_bits_size};
	wire _T_642 = _GEN_82 == a_size_lookup;
	wire _T_652 = (((_T_605 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_607;
	wire _T_654 = ~io_in_d_ready | io_in_a_ready;
	wire [159:0] a_set_wo_ready = _GEN_15[159:0];
	wire [159:0] d_clr_wo_ready = _GEN_21[159:0];
	wire _T_661 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [159:0] a_set = _GEN_16[159:0];
	wire [159:0] _inflight_T = inflight | a_set;
	wire [159:0] d_clr = _GEN_22[159:0];
	wire [159:0] _inflight_T_1 = ~d_clr;
	wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [639:0] a_opcodes_set = _GEN_19[639:0];
	wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [639:0] d_opcodes_clr = _GEN_23[639:0];
	wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [639:0] a_sizes_set = _GEN_20[639:0];
	wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_670 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [159:0] inflight_1;
	reg [639:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [639:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[639:1]};
	wire _T_696 = (io_in_d_valid & d_first_2) & _T_401;
	wire [255:0] _GEN_67 = ((d_first_done & d_first_2) & _T_401 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_68 = ((d_first_done & d_first_2) & _T_401 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire [159:0] _T_704 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_714 = _GEN_82 == c_size_lookup;
	wire [159:0] d_clr_1 = _GEN_67[159:0];
	wire [159:0] _inflight_T_4 = ~d_clr_1;
	wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0];
	wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_739 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			param <= io_in_a_bits_param;
		if (a_first_done & a_first)
			size <= io_in_a_bits_size;
		if (a_first_done & a_first)
			source <= io_in_a_bits_source;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 160'h0000000000000000000000000000000000000000;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 640'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 640'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 160'h0000000000000000000000000000000000000000;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 640'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (d_first_done)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module LevelGateway (
	clock,
	reset,
	io_interrupt,
	io_plic_valid,
	io_plic_ready,
	io_plic_complete
);
	input clock;
	input reset;
	input io_interrupt;
	output wire io_plic_valid;
	input io_plic_ready;
	input io_plic_complete;
	reg inFlight;
	wire _GEN_0 = (io_interrupt & io_plic_ready) | inFlight;
	assign io_plic_valid = io_interrupt & ~inFlight;
	always @(posedge clock)
		if (reset)
			inFlight <= 1'h0;
		else if (io_plic_complete)
			inFlight <= 1'h0;
		else
			inFlight <= _GEN_0;
endmodule
module PLICFanIn (
	io_prio_0,
	io_ip,
	io_dev,
	io_max
);
	input io_prio_0;
	input io_ip;
	output wire io_dev;
	output wire io_max;
	wire [1:0] effectivePriority_1 = {io_ip, io_prio_0};
	wire _T = 2'h2 >= effectivePriority_1;
	wire [1:0] maxPri = (_T ? 2'h2 : effectivePriority_1);
	assign io_dev = (_T ? 1'h0 : 1'h1);
	assign io_max = maxPri[0];
endmodule
module Queue_21 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_read,
	io_enq_bits_index,
	io_enq_bits_data,
	io_enq_bits_mask,
	io_enq_bits_extra_tlrr_extra_source,
	io_enq_bits_extra_tlrr_extra_size,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_read,
	io_deq_bits_index,
	io_deq_bits_data,
	io_deq_bits_mask,
	io_deq_bits_extra_tlrr_extra_source,
	io_deq_bits_extra_tlrr_extra_size
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input io_enq_bits_read;
	input [23:0] io_enq_bits_index;
	input [31:0] io_enq_bits_data;
	input [3:0] io_enq_bits_mask;
	input [7:0] io_enq_bits_extra_tlrr_extra_source;
	input [1:0] io_enq_bits_extra_tlrr_extra_size;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire io_deq_bits_read;
	output wire [23:0] io_deq_bits_index;
	output wire [31:0] io_deq_bits_data;
	output wire [3:0] io_deq_bits_mask;
	output wire [7:0] io_deq_bits_extra_tlrr_extra_source;
	output wire [1:0] io_deq_bits_extra_tlrr_extra_size;
	reg ram_read [0:0];
	wire ram_read_io_deq_bits_MPORT_en;
	wire ram_read_io_deq_bits_MPORT_addr;
	wire ram_read_io_deq_bits_MPORT_data;
	wire ram_read_MPORT_data;
	wire ram_read_MPORT_addr;
	wire ram_read_MPORT_mask;
	wire ram_read_MPORT_en;
	reg [23:0] ram_index [0:0];
	wire ram_index_io_deq_bits_MPORT_en;
	wire ram_index_io_deq_bits_MPORT_addr;
	wire [23:0] ram_index_io_deq_bits_MPORT_data;
	wire [23:0] ram_index_MPORT_data;
	wire ram_index_MPORT_addr;
	wire ram_index_MPORT_mask;
	wire ram_index_MPORT_en;
	reg [31:0] ram_data [0:0];
	wire ram_data_io_deq_bits_MPORT_en;
	wire ram_data_io_deq_bits_MPORT_addr;
	wire [31:0] ram_data_io_deq_bits_MPORT_data;
	wire [31:0] ram_data_MPORT_data;
	wire ram_data_MPORT_addr;
	wire ram_data_MPORT_mask;
	wire ram_data_MPORT_en;
	reg [3:0] ram_mask [0:0];
	wire ram_mask_io_deq_bits_MPORT_en;
	wire ram_mask_io_deq_bits_MPORT_addr;
	wire [3:0] ram_mask_io_deq_bits_MPORT_data;
	wire [3:0] ram_mask_MPORT_data;
	wire ram_mask_MPORT_addr;
	wire ram_mask_MPORT_mask;
	wire ram_mask_MPORT_en;
	reg [7:0] ram_extra_tlrr_extra_source [0:0];
	wire ram_extra_tlrr_extra_source_io_deq_bits_MPORT_en;
	wire ram_extra_tlrr_extra_source_io_deq_bits_MPORT_addr;
	wire [7:0] ram_extra_tlrr_extra_source_io_deq_bits_MPORT_data;
	wire [7:0] ram_extra_tlrr_extra_source_MPORT_data;
	wire ram_extra_tlrr_extra_source_MPORT_addr;
	wire ram_extra_tlrr_extra_source_MPORT_mask;
	wire ram_extra_tlrr_extra_source_MPORT_en;
	reg [1:0] ram_extra_tlrr_extra_size [0:0];
	wire ram_extra_tlrr_extra_size_io_deq_bits_MPORT_en;
	wire ram_extra_tlrr_extra_size_io_deq_bits_MPORT_addr;
	wire [1:0] ram_extra_tlrr_extra_size_io_deq_bits_MPORT_data;
	wire [1:0] ram_extra_tlrr_extra_size_MPORT_data;
	wire ram_extra_tlrr_extra_size_MPORT_addr;
	wire ram_extra_tlrr_extra_size_MPORT_mask;
	wire ram_extra_tlrr_extra_size_MPORT_en;
	reg maybe_full;
	wire empty = ~maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_read_io_deq_bits_MPORT_en = 1'h1;
	assign ram_read_io_deq_bits_MPORT_addr = 1'h0;
	assign ram_read_io_deq_bits_MPORT_data = ram_read[ram_read_io_deq_bits_MPORT_addr];
	assign ram_read_MPORT_data = io_enq_bits_read;
	assign ram_read_MPORT_addr = 1'h0;
	assign ram_read_MPORT_mask = 1'h1;
	assign ram_read_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_index_io_deq_bits_MPORT_en = 1'h1;
	assign ram_index_io_deq_bits_MPORT_addr = 1'h0;
	assign ram_index_io_deq_bits_MPORT_data = ram_index[ram_index_io_deq_bits_MPORT_addr];
	assign ram_index_MPORT_data = io_enq_bits_index;
	assign ram_index_MPORT_addr = 1'h0;
	assign ram_index_MPORT_mask = 1'h1;
	assign ram_index_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_data_io_deq_bits_MPORT_en = 1'h1;
	assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
	assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr];
	assign ram_data_MPORT_data = io_enq_bits_data;
	assign ram_data_MPORT_addr = 1'h0;
	assign ram_data_MPORT_mask = 1'h1;
	assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
	assign ram_mask_io_deq_bits_MPORT_addr = 1'h0;
	assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr];
	assign ram_mask_MPORT_data = io_enq_bits_mask;
	assign ram_mask_MPORT_addr = 1'h0;
	assign ram_mask_MPORT_mask = 1'h1;
	assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_extra_tlrr_extra_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_extra_tlrr_extra_source_io_deq_bits_MPORT_addr = 1'h0;
	assign ram_extra_tlrr_extra_source_io_deq_bits_MPORT_data = ram_extra_tlrr_extra_source[ram_extra_tlrr_extra_source_io_deq_bits_MPORT_addr];
	assign ram_extra_tlrr_extra_source_MPORT_data = io_enq_bits_extra_tlrr_extra_source;
	assign ram_extra_tlrr_extra_source_MPORT_addr = 1'h0;
	assign ram_extra_tlrr_extra_source_MPORT_mask = 1'h1;
	assign ram_extra_tlrr_extra_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_extra_tlrr_extra_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_extra_tlrr_extra_size_io_deq_bits_MPORT_addr = 1'h0;
	assign ram_extra_tlrr_extra_size_io_deq_bits_MPORT_data = ram_extra_tlrr_extra_size[ram_extra_tlrr_extra_size_io_deq_bits_MPORT_addr];
	assign ram_extra_tlrr_extra_size_MPORT_data = io_enq_bits_extra_tlrr_extra_size;
	assign ram_extra_tlrr_extra_size_MPORT_addr = 1'h0;
	assign ram_extra_tlrr_extra_size_MPORT_mask = 1'h1;
	assign ram_extra_tlrr_extra_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~maybe_full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_read = ram_read_io_deq_bits_MPORT_data;
	assign io_deq_bits_index = ram_index_io_deq_bits_MPORT_data;
	assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data;
	assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data;
	assign io_deq_bits_extra_tlrr_extra_source = ram_extra_tlrr_extra_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_extra_tlrr_extra_size = ram_extra_tlrr_extra_size_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_read_MPORT_en & ram_read_MPORT_mask)
			ram_read[ram_read_MPORT_addr] <= ram_read_MPORT_data;
		if (ram_index_MPORT_en & ram_index_MPORT_mask)
			ram_index[ram_index_MPORT_addr] <= ram_index_MPORT_data;
		if (ram_data_MPORT_en & ram_data_MPORT_mask)
			ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data;
		if (ram_mask_MPORT_en & ram_mask_MPORT_mask)
			ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data;
		if (ram_extra_tlrr_extra_source_MPORT_en & ram_extra_tlrr_extra_source_MPORT_mask)
			ram_extra_tlrr_extra_source[ram_extra_tlrr_extra_source_MPORT_addr] <= ram_extra_tlrr_extra_source_MPORT_data;
		if (ram_extra_tlrr_extra_size_MPORT_en & ram_extra_tlrr_extra_size_MPORT_mask)
			ram_extra_tlrr_extra_size[ram_extra_tlrr_extra_size_MPORT_addr] <= ram_extra_tlrr_extra_size_MPORT_data;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module TLPLIC (
	clock,
	reset,
	auto_int_in_0,
	auto_int_out_0,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data
);
	input clock;
	input reset;
	input auto_int_in_0;
	output wire auto_int_out_0;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [1:0] auto_in_a_bits_size;
	input [7:0] auto_in_a_bits_source;
	input [27:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_size;
	output wire [7:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [1:0] monitor_io_in_a_bits_size;
	wire [7:0] monitor_io_in_a_bits_source;
	wire [27:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_size;
	wire [7:0] monitor_io_in_d_bits_source;
	wire gateways_gateway_clock;
	wire gateways_gateway_reset;
	wire gateways_gateway_io_interrupt;
	wire gateways_gateway_io_plic_valid;
	wire gateways_gateway_io_plic_ready;
	wire gateways_gateway_io_plic_complete;
	wire fanin_io_prio_0;
	wire fanin_io_ip;
	wire fanin_io_dev;
	wire fanin_io_max;
	wire out_back_clock;
	wire out_back_reset;
	wire out_back_io_enq_ready;
	wire out_back_io_enq_valid;
	wire out_back_io_enq_bits_read;
	wire [23:0] out_back_io_enq_bits_index;
	wire [31:0] out_back_io_enq_bits_data;
	wire [3:0] out_back_io_enq_bits_mask;
	wire [7:0] out_back_io_enq_bits_extra_tlrr_extra_source;
	wire [1:0] out_back_io_enq_bits_extra_tlrr_extra_size;
	wire out_back_io_deq_ready;
	wire out_back_io_deq_valid;
	wire out_back_io_deq_bits_read;
	wire [23:0] out_back_io_deq_bits_index;
	wire [31:0] out_back_io_deq_bits_data;
	wire [3:0] out_back_io_deq_bits_mask;
	wire [7:0] out_back_io_deq_bits_extra_tlrr_extra_source;
	wire [1:0] out_back_io_deq_bits_extra_tlrr_extra_size;
	reg priority_0;
	reg threshold_0;
	reg pending_0;
	reg enables_0_0;
	wire [1:0] enableVec0_0 = {enables_0_0, 1'h0};
	reg maxDevs_0;
	reg bundleOut_0_0_REG;
	wire [2:0] out_oindex = {out_back_io_deq_bits_index[19], out_back_io_deq_bits_index[11], out_back_io_deq_bits_index[0]};
	wire [7:0] _out_backSel_T = 8'h01 << out_oindex;
	wire out_backSel_5 = _out_backSel_T[5];
	wire [23:0] out_bindex = out_back_io_deq_bits_index & 24'hf7f7fe;
	wire _out_T_3 = out_bindex == 24'h000000;
	wire out_roready_2 = (((out_back_io_deq_valid & auto_in_d_ready) & out_back_io_deq_bits_read) & out_backSel_5) & (out_bindex == 24'h000000);
	wire [7:0] _out_backMask_T_11 = (out_back_io_deq_bits_mask[3] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_9 = (out_back_io_deq_bits_mask[2] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_7 = (out_back_io_deq_bits_mask[1] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_5 = (out_back_io_deq_bits_mask[0] ? 8'hff : 8'h00);
	wire [31:0] out_backMask = {_out_backMask_T_11, _out_backMask_T_9, _out_backMask_T_7, _out_backMask_T_5};
	wire out_romask_2 = |out_backMask;
	wire out_f_roready_2 = out_roready_2 & out_romask_2;
	wire _T_5 = ~reset;
	wire claiming = out_f_roready_2 & maxDevs_0;
	wire [1:0] _claimedDevs_T = 2'h1 << claiming;
	wire claimedDevs_1 = _claimedDevs_T[1];
	wire out_woready_2 = (((out_back_io_deq_valid & auto_in_d_ready) & ~out_back_io_deq_bits_read) & out_backSel_5) & (out_bindex == 24'h000000);
	wire out_womask_2 = &out_backMask;
	wire out_f_woready_2 = out_woready_2 & out_womask_2;
	wire [31:0] _out_T_28 = out_back_io_deq_bits_data;
	wire completerDev = _out_T_28[0];
	wire [1:0] _out_completer_0_T = enableVec0_0 >> completerDev;
	wire completer_0 = out_f_woready_2 & _out_completer_0_T[0];
	wire [1:0] _completedDevs_T = 2'h1 << completerDev;
	wire [1:0] completedDevs = (completer_0 ? _completedDevs_T : 2'h0);
	wire _out_T_1 = out_bindex == 24'h000400;
	wire out_womask = &out_backMask[0];
	wire out_womask_1 = &out_backMask[1];
	wire [1:0] out_prepend = {pending_0, 1'h0};
	wire [31:0] _out_T_42 = {31'd0, maxDevs_0};
	wire out_backSel_1 = _out_backSel_T[1];
	wire out_woready_3 = (((out_back_io_deq_valid & auto_in_d_ready) & ~out_back_io_deq_bits_read) & out_backSel_1) & (out_bindex == 24'h000000);
	wire out_f_woready_3 = out_woready_3 & out_womask;
	wire out_backSel_4 = _out_backSel_T[4];
	wire out_woready_4 = (((out_back_io_deq_valid & auto_in_d_ready) & ~out_back_io_deq_bits_read) & out_backSel_4) & (out_bindex == 24'h000000);
	wire out_f_woready_4 = out_woready_4 & out_womask;
	wire [1:0] out_prepend_1 = {1'h0, threshold_0};
	wire [31:0] _out_T_73 = {30'd0, out_prepend_1};
	wire out_backSel_2 = _out_backSel_T[2];
	wire out_woready_6 = (((out_back_io_deq_valid & auto_in_d_ready) & ~out_back_io_deq_bits_read) & out_backSel_2) & (out_bindex == 24'h000000);
	wire out_f_woready_7 = out_woready_6 & out_womask_1;
	wire _GEN_37 = (3'h1 == out_oindex ? _out_T_3 : _out_T_1);
	wire _GEN_38 = (3'h2 == out_oindex ? _out_T_3 : _GEN_37);
	wire _GEN_40 = (3'h4 == out_oindex ? _out_T_3 : (3'h3 == out_oindex) | _GEN_38);
	wire _GEN_41 = (3'h5 == out_oindex ? _out_T_3 : _GEN_40);
	wire _GEN_43 = (3'h7 == out_oindex) | ((3'h6 == out_oindex) | _GEN_41);
	wire [31:0] _out_out_bits_data_WIRE_1_0 = {30'd0, out_prepend};
	wire [31:0] _out_out_bits_data_WIRE_1_1 = {31'd0, priority_0};
	wire [31:0] _GEN_45 = (3'h1 == out_oindex ? _out_out_bits_data_WIRE_1_1 : _out_out_bits_data_WIRE_1_0);
	wire [31:0] _out_out_bits_data_WIRE_1_2 = {30'd0, enableVec0_0};
	wire [31:0] _GEN_46 = (3'h2 == out_oindex ? _out_out_bits_data_WIRE_1_2 : _GEN_45);
	wire [31:0] _GEN_47 = (3'h3 == out_oindex ? 32'h00000000 : _GEN_46);
	wire [31:0] _GEN_48 = (3'h4 == out_oindex ? _out_T_73 : _GEN_47);
	wire [31:0] _GEN_49 = (3'h5 == out_oindex ? _out_T_42 : _GEN_48);
	wire [31:0] _GEN_50 = (3'h6 == out_oindex ? 32'h00000000 : _GEN_49);
	wire [31:0] _GEN_51 = (3'h7 == out_oindex ? 32'h00000000 : _GEN_50);
	wire out_bits_read = out_back_io_deq_bits_read;
	TLMonitor_34 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	LevelGateway gateways_gateway(
		.clock(gateways_gateway_clock),
		.reset(gateways_gateway_reset),
		.io_interrupt(gateways_gateway_io_interrupt),
		.io_plic_valid(gateways_gateway_io_plic_valid),
		.io_plic_ready(gateways_gateway_io_plic_ready),
		.io_plic_complete(gateways_gateway_io_plic_complete)
	);
	PLICFanIn fanin(
		.io_prio_0(fanin_io_prio_0),
		.io_ip(fanin_io_ip),
		.io_dev(fanin_io_dev),
		.io_max(fanin_io_max)
	);
	Queue_21 out_back(
		.clock(out_back_clock),
		.reset(out_back_reset),
		.io_enq_ready(out_back_io_enq_ready),
		.io_enq_valid(out_back_io_enq_valid),
		.io_enq_bits_read(out_back_io_enq_bits_read),
		.io_enq_bits_index(out_back_io_enq_bits_index),
		.io_enq_bits_data(out_back_io_enq_bits_data),
		.io_enq_bits_mask(out_back_io_enq_bits_mask),
		.io_enq_bits_extra_tlrr_extra_source(out_back_io_enq_bits_extra_tlrr_extra_source),
		.io_enq_bits_extra_tlrr_extra_size(out_back_io_enq_bits_extra_tlrr_extra_size),
		.io_deq_ready(out_back_io_deq_ready),
		.io_deq_valid(out_back_io_deq_valid),
		.io_deq_bits_read(out_back_io_deq_bits_read),
		.io_deq_bits_index(out_back_io_deq_bits_index),
		.io_deq_bits_data(out_back_io_deq_bits_data),
		.io_deq_bits_mask(out_back_io_deq_bits_mask),
		.io_deq_bits_extra_tlrr_extra_source(out_back_io_deq_bits_extra_tlrr_extra_source),
		.io_deq_bits_extra_tlrr_extra_size(out_back_io_deq_bits_extra_tlrr_extra_size)
	);
	assign auto_int_out_0 = bundleOut_0_0_REG > threshold_0;
	assign auto_in_a_ready = out_back_io_enq_ready;
	assign auto_in_d_valid = out_back_io_deq_valid;
	assign auto_in_d_bits_opcode = {2'd0, out_bits_read};
	assign auto_in_d_bits_size = out_back_io_deq_bits_extra_tlrr_extra_size;
	assign auto_in_d_bits_source = out_back_io_deq_bits_extra_tlrr_extra_source;
	assign auto_in_d_bits_data = (_GEN_43 ? _GEN_51 : 32'h00000000);
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = out_back_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = out_back_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = {2'd0, out_bits_read};
	assign monitor_io_in_d_bits_size = out_back_io_deq_bits_extra_tlrr_extra_size;
	assign monitor_io_in_d_bits_source = out_back_io_deq_bits_extra_tlrr_extra_source;
	assign gateways_gateway_clock = clock;
	assign gateways_gateway_reset = reset;
	assign gateways_gateway_io_interrupt = auto_int_in_0;
	assign gateways_gateway_io_plic_ready = ~pending_0;
	assign gateways_gateway_io_plic_complete = completedDevs[1];
	assign fanin_io_prio_0 = priority_0;
	assign fanin_io_ip = enables_0_0 & pending_0;
	assign out_back_clock = clock;
	assign out_back_reset = reset;
	assign out_back_io_enq_valid = auto_in_a_valid;
	assign out_back_io_enq_bits_read = auto_in_a_bits_opcode == 3'h4;
	assign out_back_io_enq_bits_index = auto_in_a_bits_address[25:2];
	assign out_back_io_enq_bits_data = auto_in_a_bits_data;
	assign out_back_io_enq_bits_mask = auto_in_a_bits_mask;
	assign out_back_io_enq_bits_extra_tlrr_extra_source = auto_in_a_bits_source;
	assign out_back_io_enq_bits_extra_tlrr_extra_size = auto_in_a_bits_size;
	assign out_back_io_deq_ready = auto_in_d_ready;
	always @(posedge clock) begin
		if (out_f_woready_3)
			priority_0 <= out_back_io_deq_bits_data[0];
		if (out_f_woready_4)
			threshold_0 <= out_back_io_deq_bits_data[0];
		if (reset)
			pending_0 <= 1'h0;
		else if (claimedDevs_1 | gateways_gateway_io_plic_valid)
			pending_0 <= ~claimedDevs_1;
		if (out_f_woready_7)
			enables_0_0 <= out_back_io_deq_bits_data[1];
		maxDevs_0 <= fanin_io_dev;
		bundleOut_0_0_REG <= fanin_io_max;
	end
endmodule
module ClockSinkDomain (
	auto_plic_int_in_0,
	auto_plic_int_out_0,
	auto_plic_in_a_ready,
	auto_plic_in_a_valid,
	auto_plic_in_a_bits_opcode,
	auto_plic_in_a_bits_param,
	auto_plic_in_a_bits_size,
	auto_plic_in_a_bits_source,
	auto_plic_in_a_bits_address,
	auto_plic_in_a_bits_mask,
	auto_plic_in_a_bits_data,
	auto_plic_in_a_bits_corrupt,
	auto_plic_in_d_ready,
	auto_plic_in_d_valid,
	auto_plic_in_d_bits_opcode,
	auto_plic_in_d_bits_size,
	auto_plic_in_d_bits_source,
	auto_plic_in_d_bits_data,
	auto_clock_in_clock,
	auto_clock_in_reset
);
	input auto_plic_int_in_0;
	output wire auto_plic_int_out_0;
	output wire auto_plic_in_a_ready;
	input auto_plic_in_a_valid;
	input [2:0] auto_plic_in_a_bits_opcode;
	input [2:0] auto_plic_in_a_bits_param;
	input [1:0] auto_plic_in_a_bits_size;
	input [7:0] auto_plic_in_a_bits_source;
	input [27:0] auto_plic_in_a_bits_address;
	input [3:0] auto_plic_in_a_bits_mask;
	input [31:0] auto_plic_in_a_bits_data;
	input auto_plic_in_a_bits_corrupt;
	input auto_plic_in_d_ready;
	output wire auto_plic_in_d_valid;
	output wire [2:0] auto_plic_in_d_bits_opcode;
	output wire [1:0] auto_plic_in_d_bits_size;
	output wire [7:0] auto_plic_in_d_bits_source;
	output wire [31:0] auto_plic_in_d_bits_data;
	input auto_clock_in_clock;
	input auto_clock_in_reset;
	wire plic_clock;
	wire plic_reset;
	wire plic_auto_int_in_0;
	wire plic_auto_int_out_0;
	wire plic_auto_in_a_ready;
	wire plic_auto_in_a_valid;
	wire [2:0] plic_auto_in_a_bits_opcode;
	wire [2:0] plic_auto_in_a_bits_param;
	wire [1:0] plic_auto_in_a_bits_size;
	wire [7:0] plic_auto_in_a_bits_source;
	wire [27:0] plic_auto_in_a_bits_address;
	wire [3:0] plic_auto_in_a_bits_mask;
	wire [31:0] plic_auto_in_a_bits_data;
	wire plic_auto_in_a_bits_corrupt;
	wire plic_auto_in_d_ready;
	wire plic_auto_in_d_valid;
	wire [2:0] plic_auto_in_d_bits_opcode;
	wire [1:0] plic_auto_in_d_bits_size;
	wire [7:0] plic_auto_in_d_bits_source;
	wire [31:0] plic_auto_in_d_bits_data;
	TLPLIC plic(
		.clock(plic_clock),
		.reset(plic_reset),
		.auto_int_in_0(plic_auto_int_in_0),
		.auto_int_out_0(plic_auto_int_out_0),
		.auto_in_a_ready(plic_auto_in_a_ready),
		.auto_in_a_valid(plic_auto_in_a_valid),
		.auto_in_a_bits_opcode(plic_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(plic_auto_in_a_bits_param),
		.auto_in_a_bits_size(plic_auto_in_a_bits_size),
		.auto_in_a_bits_source(plic_auto_in_a_bits_source),
		.auto_in_a_bits_address(plic_auto_in_a_bits_address),
		.auto_in_a_bits_mask(plic_auto_in_a_bits_mask),
		.auto_in_a_bits_data(plic_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(plic_auto_in_a_bits_corrupt),
		.auto_in_d_ready(plic_auto_in_d_ready),
		.auto_in_d_valid(plic_auto_in_d_valid),
		.auto_in_d_bits_opcode(plic_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(plic_auto_in_d_bits_size),
		.auto_in_d_bits_source(plic_auto_in_d_bits_source),
		.auto_in_d_bits_data(plic_auto_in_d_bits_data)
	);
	assign auto_plic_int_out_0 = plic_auto_int_out_0;
	assign auto_plic_in_a_ready = plic_auto_in_a_ready;
	assign auto_plic_in_d_valid = plic_auto_in_d_valid;
	assign auto_plic_in_d_bits_opcode = plic_auto_in_d_bits_opcode;
	assign auto_plic_in_d_bits_size = plic_auto_in_d_bits_size;
	assign auto_plic_in_d_bits_source = plic_auto_in_d_bits_source;
	assign auto_plic_in_d_bits_data = plic_auto_in_d_bits_data;
	assign plic_clock = auto_clock_in_clock;
	assign plic_reset = auto_clock_in_reset;
	assign plic_auto_int_in_0 = auto_plic_int_in_0;
	assign plic_auto_in_a_valid = auto_plic_in_a_valid;
	assign plic_auto_in_a_bits_opcode = auto_plic_in_a_bits_opcode;
	assign plic_auto_in_a_bits_param = auto_plic_in_a_bits_param;
	assign plic_auto_in_a_bits_size = auto_plic_in_a_bits_size;
	assign plic_auto_in_a_bits_source = auto_plic_in_a_bits_source;
	assign plic_auto_in_a_bits_address = auto_plic_in_a_bits_address;
	assign plic_auto_in_a_bits_mask = auto_plic_in_a_bits_mask;
	assign plic_auto_in_a_bits_data = auto_plic_in_a_bits_data;
	assign plic_auto_in_a_bits_corrupt = auto_plic_in_a_bits_corrupt;
	assign plic_auto_in_d_ready = auto_plic_in_d_ready;
endmodule
module TLMonitor_35 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [1:0] io_in_a_bits_size;
	input [7:0] io_in_a_bits_source;
	input [25:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_size;
	input [7:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_4 = io_in_a_bits_source <= 8'h9f;
	wire [4:0] _is_aligned_mask_T_1 = 5'h03 << io_in_a_bits_size;
	wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0];
	wire [25:0] _GEN_71 = {24'd0, is_aligned_mask};
	wire [25:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 26'h0000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 2'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_10 = ~_source_ok_T_4;
	wire _T_20 = io_in_a_bits_opcode == 3'h6;
	wire [25:0] _T_33 = io_in_a_bits_address ^ 26'h2000000;
	wire [26:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [26:0] _T_36 = $signed(_T_34) & -27'sh0010000;
	wire _T_37 = $signed(_T_36) == 27'sh0000000;
	wire _T_69 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_73 = ~io_in_a_bits_mask;
	wire _T_74 = _T_73 == 4'h0;
	wire _T_78 = ~io_in_a_bits_corrupt;
	wire _T_82 = io_in_a_bits_opcode == 3'h7;
	wire _T_135 = io_in_a_bits_param != 3'h0;
	wire _T_148 = io_in_a_bits_opcode == 3'h4;
	wire _T_164 = io_in_a_bits_size <= 2'h2;
	wire _T_172 = _T_164 & _T_37;
	wire _T_183 = io_in_a_bits_param == 3'h0;
	wire _T_187 = io_in_a_bits_mask == mask;
	wire _T_195 = io_in_a_bits_opcode == 3'h0;
	wire _T_218 = _source_ok_T_4 & _T_172;
	wire _T_236 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_273 = ~mask;
	wire [3:0] _T_274 = io_in_a_bits_mask & _T_273;
	wire _T_275 = _T_274 == 4'h0;
	wire _T_279 = io_in_a_bits_opcode == 3'h2;
	wire _T_309 = io_in_a_bits_param <= 3'h4;
	wire _T_317 = io_in_a_bits_opcode == 3'h3;
	wire _T_347 = io_in_a_bits_param <= 3'h3;
	wire _T_355 = io_in_a_bits_opcode == 3'h5;
	wire _T_385 = io_in_a_bits_param <= 3'h1;
	wire _T_397 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_10 = io_in_d_bits_source <= 8'h9f;
	wire _T_401 = io_in_d_bits_opcode == 3'h6;
	wire _T_405 = io_in_d_bits_size >= 2'h2;
	wire _T_421 = io_in_d_bits_opcode == 3'h4;
	wire _T_449 = io_in_d_bits_opcode == 3'h5;
	wire _T_478 = io_in_d_bits_opcode == 3'h0;
	wire _T_495 = io_in_d_bits_opcode == 3'h1;
	wire _T_513 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [1:0] size;
	reg [7:0] source;
	reg [25:0] address;
	wire _T_543 = io_in_a_valid & ~a_first;
	wire _T_544 = io_in_a_bits_opcode == opcode;
	wire _T_548 = io_in_a_bits_param == param;
	wire _T_552 = io_in_a_bits_size == size;
	wire _T_556 = io_in_a_bits_source == source;
	wire _T_560 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] size_1;
	reg [7:0] source_1;
	wire _T_567 = io_in_d_valid & ~d_first;
	wire _T_568 = io_in_d_bits_opcode == opcode_1;
	wire _T_576 = io_in_d_bits_size == size_1;
	wire _T_580 = io_in_d_bits_source == source_1;
	reg [159:0] inflight;
	reg [639:0] inflight_opcodes;
	reg [639:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [10:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [639:0] _GEN_73 = {624'd0, _a_opcode_lookup_T_5};
	wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [639:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[639:1]};
	wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [639:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[639:1]};
	wire _T_594 = io_in_a_valid & a_first_1;
	wire [255:0] _a_set_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_a_bits_source;
	wire _T_597 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1;
	wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [10:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [2050:0] _GEN_1 = {2047'd0, a_opcodes_set_interm};
	wire [2050:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? _a_sizes_set_interm_T_1 : 3'h0);
	wire [2049:0] _GEN_2 = {2047'd0, a_sizes_set_interm};
	wire [2049:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [159:0] _T_599 = inflight >> io_in_a_bits_source;
	wire _T_601 = ~_T_599[0];
	wire [255:0] _GEN_16 = (a_first_done & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2050:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 2051'h0);
	wire [2049:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 2050'h0);
	wire _T_605 = io_in_d_valid & d_first_1;
	wire _T_607 = ~_T_401;
	wire _T_608 = (io_in_d_valid & d_first_1) & ~_T_401;
	wire [255:0] _d_clr_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_d_bits_source;
	wire [2062:0] _GEN_3 = {2047'd0, _a_opcode_lookup_T_5};
	wire [2062:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [255:0] _GEN_22 = ((d_first_done & d_first_1) & _T_607 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_23 = ((d_first_done & d_first_1) & _T_607 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_594 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [159:0] _T_618 = inflight >> io_in_d_bits_source;
	wire _T_620 = _T_618[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_625 = io_in_d_bits_opcode == _GEN_40;
	wire _T_626 = (io_in_d_bits_opcode == _GEN_32) | _T_625;
	wire _T_630 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_637 = io_in_d_bits_opcode == _GEN_56;
	wire _T_638 = (io_in_d_bits_opcode == _GEN_48) | _T_637;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {2'd0, io_in_d_bits_size};
	wire _T_642 = _GEN_82 == a_size_lookup;
	wire _T_652 = (((_T_605 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_607;
	wire _T_654 = ~io_in_d_ready | io_in_a_ready;
	wire [159:0] a_set = _GEN_16[159:0];
	wire [159:0] _inflight_T = inflight | a_set;
	wire [159:0] d_clr = _GEN_22[159:0];
	wire [159:0] _inflight_T_1 = ~d_clr;
	wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [639:0] a_opcodes_set = _GEN_19[639:0];
	wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [639:0] d_opcodes_clr = _GEN_23[639:0];
	wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [639:0] a_sizes_set = _GEN_20[639:0];
	wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_663 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [159:0] inflight_1;
	reg [639:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [639:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[639:1]};
	wire _T_689 = (io_in_d_valid & d_first_2) & _T_401;
	wire [255:0] _GEN_67 = ((d_first_done & d_first_2) & _T_401 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_68 = ((d_first_done & d_first_2) & _T_401 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire [159:0] _T_697 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_707 = _GEN_82 == c_size_lookup;
	wire [159:0] d_clr_1 = _GEN_67[159:0];
	wire [159:0] _inflight_T_4 = ~d_clr_1;
	wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0];
	wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_727 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			param <= io_in_a_bits_param;
		if (a_first_done & a_first)
			size <= io_in_a_bits_size;
		if (a_first_done & a_first)
			source <= io_in_a_bits_source;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 160'h0000000000000000000000000000000000000000;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 640'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 640'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 160'h0000000000000000000000000000000000000000;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 640'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (d_first_done)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module CLINT (
	clock,
	reset,
	auto_int_out_0,
	auto_int_out_1,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	io_rtcTick
);
	input clock;
	input reset;
	output wire auto_int_out_0;
	output wire auto_int_out_1;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [1:0] auto_in_a_bits_size;
	input [7:0] auto_in_a_bits_source;
	input [25:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_size;
	output wire [7:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input io_rtcTick;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [1:0] monitor_io_in_a_bits_size;
	wire [7:0] monitor_io_in_a_bits_source;
	wire [25:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_size;
	wire [7:0] monitor_io_in_d_bits_source;
	reg [63:0] time_;
	wire [63:0] _time_T_1 = time_ + 64'h0000000000000001;
	reg [63:0] timecmp_0;
	reg ipi_0;
	wire [7:0] oldBytes__0 = timecmp_0[7:0];
	wire [7:0] oldBytes__1 = timecmp_0[15:8];
	wire [7:0] oldBytes__2 = timecmp_0[23:16];
	wire [7:0] oldBytes__3 = timecmp_0[31:24];
	wire [7:0] oldBytes__4 = timecmp_0[39:32];
	wire [7:0] oldBytes__5 = timecmp_0[47:40];
	wire [7:0] oldBytes__6 = timecmp_0[55:48];
	wire [7:0] oldBytes__7 = timecmp_0[63:56];
	wire in_bits_read = auto_in_a_bits_opcode == 3'h4;
	wire [13:0] in_bits_index = auto_in_a_bits_address[15:2];
	wire [2:0] out_iindex = {in_bits_index[13], in_bits_index[12], in_bits_index[0]};
	wire [13:0] out_findex = in_bits_index & 14'h0ffe;
	wire _out_T_6 = out_findex == 14'h0ffe;
	wire _out_T_2 = out_findex == 14'h0000;
	wire [7:0] _out_backSel_T = 8'h01 << out_iindex;
	wire out_backSel_2 = _out_backSel_T[2];
	wire out_woready_14 = (((auto_in_a_valid & auto_in_d_ready) & ~in_bits_read) & out_backSel_2) & (out_findex == 14'h0000);
	wire [7:0] _out_backMask_T_11 = (auto_in_a_bits_mask[3] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_9 = (auto_in_a_bits_mask[2] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_7 = (auto_in_a_bits_mask[1] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_5 = (auto_in_a_bits_mask[0] ? 8'hff : 8'h00);
	wire [31:0] out_backMask = {_out_backMask_T_11, _out_backMask_T_9, _out_backMask_T_7, _out_backMask_T_5};
	wire out_womask_14 = &out_backMask[7:0];
	wire out_f_woready_14 = out_woready_14 & out_womask_14;
	wire out_womask_15 = &out_backMask[15:8];
	wire out_f_woready_15 = out_woready_14 & out_womask_15;
	wire out_womask_16 = &out_backMask[23:16];
	wire out_f_woready_16 = out_woready_14 & out_womask_16;
	wire out_womask_17 = &out_backMask[31:24];
	wire out_f_woready_17 = out_woready_14 & out_womask_17;
	wire out_backSel_3 = _out_backSel_T[3];
	wire out_woready_2 = (((auto_in_a_valid & auto_in_d_ready) & ~in_bits_read) & out_backSel_3) & (out_findex == 14'h0000);
	wire out_f_woready_2 = out_woready_2 & out_womask_14;
	wire out_f_woready_3 = out_woready_2 & out_womask_15;
	wire out_f_woready_4 = out_woready_2 & out_womask_16;
	wire out_f_woready_5 = out_woready_2 & out_womask_17;
	wire [7:0] newBytes__1 = (out_f_woready_15 ? auto_in_a_bits_data[15:8] : oldBytes__1);
	wire [7:0] newBytes__0 = (out_f_woready_14 ? auto_in_a_bits_data[7:0] : oldBytes__0);
	wire [7:0] newBytes__3 = (out_f_woready_17 ? auto_in_a_bits_data[31:24] : oldBytes__3);
	wire [7:0] newBytes__2 = (out_f_woready_16 ? auto_in_a_bits_data[23:16] : oldBytes__2);
	wire [7:0] newBytes__5 = (out_f_woready_3 ? auto_in_a_bits_data[15:8] : oldBytes__5);
	wire [7:0] newBytes__4 = (out_f_woready_2 ? auto_in_a_bits_data[7:0] : oldBytes__4);
	wire [7:0] newBytes__7 = (out_f_woready_5 ? auto_in_a_bits_data[31:24] : oldBytes__7);
	wire [7:0] newBytes__6 = (out_f_woready_4 ? auto_in_a_bits_data[23:16] : oldBytes__6);
	wire [63:0] _timecmp_0_T = {newBytes__7, newBytes__6, newBytes__5, newBytes__4, newBytes__3, newBytes__2, newBytes__1, newBytes__0};
	wire [7:0] oldBytes_1_0 = time_[7:0];
	wire [7:0] oldBytes_1_1 = time_[15:8];
	wire [7:0] oldBytes_1_2 = time_[23:16];
	wire [7:0] oldBytes_1_3 = time_[31:24];
	wire [7:0] oldBytes_1_4 = time_[39:32];
	wire [7:0] oldBytes_1_5 = time_[47:40];
	wire [7:0] oldBytes_1_6 = time_[55:48];
	wire [7:0] oldBytes_1_7 = time_[63:56];
	wire out_backSel_4 = _out_backSel_T[4];
	wire out_woready_6 = (((auto_in_a_valid & auto_in_d_ready) & ~in_bits_read) & out_backSel_4) & (out_findex == 14'h0ffe);
	wire out_f_woready_6 = out_woready_6 & out_womask_14;
	wire out_f_woready_7 = out_woready_6 & out_womask_15;
	wire out_f_woready_8 = out_woready_6 & out_womask_16;
	wire out_f_woready_9 = out_woready_6 & out_womask_17;
	wire out_backSel_5 = _out_backSel_T[5];
	wire out_woready_10 = (((auto_in_a_valid & auto_in_d_ready) & ~in_bits_read) & out_backSel_5) & (out_findex == 14'h0ffe);
	wire out_f_woready_10 = out_woready_10 & out_womask_14;
	wire out_f_woready_11 = out_woready_10 & out_womask_15;
	wire out_f_woready_12 = out_woready_10 & out_womask_16;
	wire out_f_woready_13 = out_woready_10 & out_womask_17;
	wire [7:0] newBytes_1_1 = (out_f_woready_7 ? auto_in_a_bits_data[15:8] : oldBytes_1_1);
	wire [7:0] newBytes_1_0 = (out_f_woready_6 ? auto_in_a_bits_data[7:0] : oldBytes_1_0);
	wire [7:0] newBytes_1_3 = (out_f_woready_9 ? auto_in_a_bits_data[31:24] : oldBytes_1_3);
	wire [7:0] newBytes_1_2 = (out_f_woready_8 ? auto_in_a_bits_data[23:16] : oldBytes_1_2);
	wire [7:0] newBytes_1_5 = (out_f_woready_11 ? auto_in_a_bits_data[15:8] : oldBytes_1_5);
	wire [7:0] newBytes_1_4 = (out_f_woready_10 ? auto_in_a_bits_data[7:0] : oldBytes_1_4);
	wire [7:0] newBytes_1_7 = (out_f_woready_13 ? auto_in_a_bits_data[31:24] : oldBytes_1_7);
	wire [7:0] newBytes_1_6 = (out_f_woready_12 ? auto_in_a_bits_data[23:16] : oldBytes_1_6);
	wire [63:0] _time_T_2 = {newBytes_1_7, newBytes_1_6, newBytes_1_5, newBytes_1_4, newBytes_1_3, newBytes_1_2, newBytes_1_1, newBytes_1_0};
	wire out_wimask = &out_backMask[0];
	wire out_frontSel_0 = _out_backSel_T[0];
	wire out_wivalid_0 = (((auto_in_a_valid & auto_in_d_ready) & ~in_bits_read) & out_frontSel_0) & (out_findex == 14'h0000);
	wire out_f_wivalid = out_wivalid_0 & out_wimask;
	wire [1:0] out_prepend = {1'h0, ipi_0};
	wire [31:0] _out_T_28 = {30'd0, out_prepend};
	wire [31:0] out_prepend_3 = {oldBytes__7, oldBytes__6, oldBytes__5, oldBytes__4};
	wire [31:0] out_prepend_6 = {oldBytes_1_3, oldBytes_1_2, oldBytes_1_1, oldBytes_1_0};
	wire [31:0] out_prepend_9 = {oldBytes_1_7, oldBytes_1_6, oldBytes_1_5, oldBytes_1_4};
	wire [31:0] out_prepend_12 = {oldBytes__3, oldBytes__2, oldBytes__1, oldBytes__0};
	wire _GEN_54 = (3'h2 == out_iindex ? _out_T_2 : (3'h1 == out_iindex) | _out_T_2);
	wire _GEN_55 = (3'h3 == out_iindex ? _out_T_2 : _GEN_54);
	wire _GEN_56 = (3'h4 == out_iindex ? _out_T_6 : _GEN_55);
	wire _GEN_57 = (3'h5 == out_iindex ? _out_T_6 : _GEN_56);
	wire _GEN_59 = (3'h7 == out_iindex) | ((3'h6 == out_iindex) | _GEN_57);
	wire [31:0] _GEN_61 = (3'h1 == out_iindex ? 32'h00000000 : _out_T_28);
	wire [31:0] _GEN_62 = (3'h2 == out_iindex ? out_prepend_12 : _GEN_61);
	wire [31:0] _GEN_63 = (3'h3 == out_iindex ? out_prepend_3 : _GEN_62);
	wire [31:0] _GEN_64 = (3'h4 == out_iindex ? out_prepend_6 : _GEN_63);
	wire [31:0] _GEN_65 = (3'h5 == out_iindex ? out_prepend_9 : _GEN_64);
	wire [31:0] _GEN_66 = (3'h6 == out_iindex ? 32'h00000000 : _GEN_65);
	wire [31:0] _GEN_67 = (3'h7 == out_iindex ? 32'h00000000 : _GEN_66);
	TLMonitor_35 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	assign auto_int_out_0 = ipi_0;
	assign auto_int_out_1 = time_ >= timecmp_0;
	assign auto_in_a_ready = auto_in_d_ready;
	assign auto_in_d_valid = auto_in_a_valid;
	assign auto_in_d_bits_opcode = {2'd0, in_bits_read};
	assign auto_in_d_bits_size = auto_in_a_bits_size;
	assign auto_in_d_bits_source = auto_in_a_bits_source;
	assign auto_in_d_bits_data = (_GEN_59 ? _GEN_67 : 32'h00000000);
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_in_d_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_in_a_valid;
	assign monitor_io_in_d_bits_opcode = {2'd0, in_bits_read};
	assign monitor_io_in_d_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_d_bits_source = auto_in_a_bits_source;
	always @(posedge clock) begin
		if (reset)
			time_ <= 64'h0000000000000000;
		else if (((((((out_f_woready_6 | out_f_woready_7) | out_f_woready_8) | out_f_woready_9) | out_f_woready_10) | out_f_woready_11) | out_f_woready_12) | out_f_woready_13)
			time_ <= _time_T_2;
		else if (io_rtcTick)
			time_ <= _time_T_1;
		if (((((((out_f_woready_14 | out_f_woready_15) | out_f_woready_16) | out_f_woready_17) | out_f_woready_2) | out_f_woready_3) | out_f_woready_4) | out_f_woready_5)
			timecmp_0 <= _timecmp_0_T;
		if (reset)
			ipi_0 <= 1'h0;
		else if (out_f_wivalid)
			ipi_0 <= auto_in_a_bits_data[0];
	end
endmodule
module TLMonitor_36 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_address,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [8:0] io_in_a_bits_address;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [1:0] io_in_d_bits_size;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire [8:0] _is_aligned_T = io_in_a_bits_address & 9'h003;
	wire is_aligned = _is_aligned_T == 9'h000;
	wire [9:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_15 = io_in_a_bits_opcode == 3'h6;
	wire [9:0] _T_23 = $signed(_T_7) & 10'sh200;
	wire _T_24 = $signed(_T_23) == 10'sh000;
	wire _T_69 = io_in_a_bits_opcode == 3'h7;
	wire _T_127 = io_in_a_bits_opcode == 3'h4;
	wire _T_167 = io_in_a_bits_opcode == 3'h0;
	wire _T_201 = io_in_a_bits_opcode == 3'h1;
	wire _T_236 = io_in_a_bits_opcode == 3'h2;
	wire _T_266 = io_in_a_bits_opcode == 3'h3;
	wire _T_296 = io_in_a_bits_opcode == 3'h5;
	wire _T_330 = io_in_d_bits_opcode <= 3'h6;
	wire _T_334 = io_in_d_bits_opcode == 3'h6;
	wire _T_338 = io_in_d_bits_size >= 2'h2;
	wire _T_342 = io_in_d_bits_param == 2'h0;
	wire _T_346 = ~io_in_d_bits_corrupt;
	wire _T_350 = ~io_in_d_bits_denied;
	wire _T_354 = io_in_d_bits_opcode == 3'h4;
	wire _T_365 = io_in_d_bits_param <= 2'h2;
	wire _T_369 = io_in_d_bits_param != 2'h2;
	wire _T_382 = io_in_d_bits_opcode == 3'h5;
	wire _T_402 = _T_350 | io_in_d_bits_corrupt;
	wire _T_411 = io_in_d_bits_opcode == 3'h0;
	wire _T_428 = io_in_d_bits_opcode == 3'h1;
	wire _T_446 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [8:0] address;
	wire _T_476 = io_in_a_valid & ~a_first;
	wire _T_477 = io_in_a_bits_opcode == opcode;
	wire _T_493 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [1:0] size_1;
	reg sink;
	reg denied;
	wire _T_500 = io_in_d_valid & ~d_first;
	wire _T_501 = io_in_d_bits_opcode == opcode_1;
	wire _T_505 = io_in_d_bits_param == param_1;
	wire _T_509 = io_in_d_bits_size == size_1;
	wire _T_517 = io_in_d_bits_sink == sink;
	wire _T_521 = io_in_d_bits_denied == denied;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [3:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_71 = {12'd0, inflight_opcodes};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_71 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [15:0] _GEN_73 = {12'd0, inflight_sizes};
	wire [15:0] _a_size_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_527 = io_in_a_valid & a_first_1;
	wire _T_530 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _a_opcodes_set_T_1 = {15'd0, a_opcodes_set_interm};
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? 3'h5 : 3'h0);
	wire [17:0] _a_sizes_set_T_1 = {15'd0, a_sizes_set_interm};
	wire _T_534 = ~inflight;
	wire [1:0] _GEN_16 = (a_first_done & a_first_1 ? 2'h1 : 2'h0);
	wire [18:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [17:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 18'h00000);
	wire _T_538 = io_in_d_valid & d_first_1;
	wire _T_540 = ~_T_334;
	wire _T_541 = (io_in_d_valid & d_first_1) & ~_T_334;
	wire [30:0] _d_opcodes_clr_T_5 = {15'd0, _a_opcode_lookup_T_5};
	wire [1:0] _GEN_22 = ((d_first_done & d_first_1) & _T_540 ? 2'h1 : 2'h0);
	wire [30:0] _GEN_23 = ((d_first_done & d_first_1) & _T_540 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire _T_553 = inflight | _T_527;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_558 = io_in_d_bits_opcode == _GEN_40;
	wire _T_559 = (io_in_d_bits_opcode == _GEN_32) | _T_558;
	wire _T_563 = 2'h2 == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_570 = io_in_d_bits_opcode == _GEN_56;
	wire _T_571 = (io_in_d_bits_opcode == _GEN_48) | _T_570;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_75 = {2'd0, io_in_d_bits_size};
	wire _T_575 = _GEN_75 == a_size_lookup;
	wire _T_585 = ((_T_538 & a_first_1) & io_in_a_valid) & _T_540;
	wire _T_587 = ~io_in_d_ready | io_in_a_ready;
	wire a_set = _GEN_16[0];
	wire d_clr = _GEN_22[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [3:0] a_sizes_set = _GEN_20[3:0];
	wire [3:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [3:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_596 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [3:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [15:0] _GEN_78 = {12'd0, inflight_sizes_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_78 & _a_opcode_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_622 = (io_in_d_valid & d_first_2) & _T_334;
	wire [30:0] _GEN_68 = ((d_first_done & d_first_2) & _T_334 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_640 = _GEN_75 == c_size_lookup;
	wire [3:0] d_opcodes_clr_1 = _GEN_68[3:0];
	wire [3:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [3:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			param_1 <= io_in_d_bits_param;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			sink <= io_in_d_bits_sink;
		if (d_first_done & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 4'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 4'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module TLXbar_8 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_address,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_1_a_ready,
	auto_out_1_a_valid,
	auto_out_1_a_bits_opcode,
	auto_out_1_a_bits_address,
	auto_out_1_a_bits_data,
	auto_out_1_d_ready,
	auto_out_1_d_valid,
	auto_out_1_d_bits_opcode,
	auto_out_1_d_bits_data,
	auto_out_0_a_ready,
	auto_out_0_a_valid,
	auto_out_0_a_bits_opcode,
	auto_out_0_a_bits_address,
	auto_out_0_a_bits_data,
	auto_out_0_d_ready,
	auto_out_0_d_valid,
	auto_out_0_d_bits_opcode,
	auto_out_0_d_bits_param,
	auto_out_0_d_bits_size,
	auto_out_0_d_bits_sink,
	auto_out_0_d_bits_denied,
	auto_out_0_d_bits_data,
	auto_out_0_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [8:0] auto_in_a_bits_address;
	input [31:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_1_a_ready;
	output wire auto_out_1_a_valid;
	output wire [2:0] auto_out_1_a_bits_opcode;
	output wire [6:0] auto_out_1_a_bits_address;
	output wire [31:0] auto_out_1_a_bits_data;
	output wire auto_out_1_d_ready;
	input auto_out_1_d_valid;
	input [2:0] auto_out_1_d_bits_opcode;
	input [31:0] auto_out_1_d_bits_data;
	input auto_out_0_a_ready;
	output wire auto_out_0_a_valid;
	output wire [2:0] auto_out_0_a_bits_opcode;
	output wire [8:0] auto_out_0_a_bits_address;
	output wire [31:0] auto_out_0_a_bits_data;
	output wire auto_out_0_d_ready;
	input auto_out_0_d_valid;
	input [2:0] auto_out_0_d_bits_opcode;
	input [1:0] auto_out_0_d_bits_param;
	input [1:0] auto_out_0_d_bits_size;
	input auto_out_0_d_bits_sink;
	input auto_out_0_d_bits_denied;
	input [31:0] auto_out_0_d_bits_data;
	input auto_out_0_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [8:0] monitor_io_in_a_bits_address;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [1:0] monitor_io_in_d_bits_size;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire [9:0] _requestAIO_T_1 = {1'b0, $signed(auto_in_a_bits_address)};
	wire [9:0] _requestAIO_T_3 = $signed(_requestAIO_T_1) & 10'sh1c0;
	wire _requestAIO_T_4 = $signed(_requestAIO_T_3) == 10'sh000;
	wire [8:0] _requestAIO_T_5 = auto_in_a_bits_address ^ 9'h044;
	wire [9:0] _requestAIO_T_6 = {1'b0, $signed(_requestAIO_T_5)};
	wire [9:0] _requestAIO_T_8 = $signed(_requestAIO_T_6) & 10'sh1f4;
	wire _requestAIO_T_9 = $signed(_requestAIO_T_8) == 10'sh000;
	wire [8:0] _requestAIO_T_10 = auto_in_a_bits_address ^ 9'h058;
	wire [9:0] _requestAIO_T_11 = {1'b0, $signed(_requestAIO_T_10)};
	wire [9:0] _requestAIO_T_13 = $signed(_requestAIO_T_11) & 10'sh1f8;
	wire _requestAIO_T_14 = $signed(_requestAIO_T_13) == 10'sh000;
	wire [8:0] _requestAIO_T_15 = auto_in_a_bits_address ^ 9'h060;
	wire [9:0] _requestAIO_T_16 = {1'b0, $signed(_requestAIO_T_15)};
	wire [9:0] _requestAIO_T_18 = $signed(_requestAIO_T_16) & 10'sh1e0;
	wire _requestAIO_T_19 = $signed(_requestAIO_T_18) == 10'sh000;
	wire [8:0] _requestAIO_T_20 = auto_in_a_bits_address ^ 9'h080;
	wire [9:0] _requestAIO_T_21 = {1'b0, $signed(_requestAIO_T_20)};
	wire [9:0] _requestAIO_T_23 = $signed(_requestAIO_T_21) & 10'sh180;
	wire _requestAIO_T_24 = $signed(_requestAIO_T_23) == 10'sh000;
	wire [8:0] _requestAIO_T_25 = auto_in_a_bits_address ^ 9'h100;
	wire [9:0] _requestAIO_T_26 = {1'b0, $signed(_requestAIO_T_25)};
	wire [9:0] _requestAIO_T_28 = $signed(_requestAIO_T_26) & 10'sh100;
	wire _requestAIO_T_29 = $signed(_requestAIO_T_28) == 10'sh000;
	wire requestAIO_0_0 = ((((_requestAIO_T_4 | _requestAIO_T_9) | _requestAIO_T_14) | _requestAIO_T_19) | _requestAIO_T_24) | _requestAIO_T_29;
	wire [8:0] _requestAIO_T_35 = auto_in_a_bits_address ^ 9'h040;
	wire [9:0] _requestAIO_T_36 = {1'b0, $signed(_requestAIO_T_35)};
	wire [9:0] _requestAIO_T_38 = $signed(_requestAIO_T_36) & 10'sh1f4;
	wire _requestAIO_T_39 = $signed(_requestAIO_T_38) == 10'sh000;
	wire [8:0] _requestAIO_T_40 = auto_in_a_bits_address ^ 9'h050;
	wire [9:0] _requestAIO_T_41 = {1'b0, $signed(_requestAIO_T_40)};
	wire [9:0] _requestAIO_T_43 = $signed(_requestAIO_T_41) & 10'sh1f8;
	wire _requestAIO_T_44 = $signed(_requestAIO_T_43) == 10'sh000;
	wire requestAIO_0_1 = _requestAIO_T_39 | _requestAIO_T_44;
	reg beatsLeft;
	wire idle = ~beatsLeft;
	wire latch = idle & auto_in_d_ready;
	wire [1:0] readys_valid = {auto_out_1_d_valid, auto_out_0_d_valid};
	wire _readys_T_3 = ~reset;
	reg [1:0] readys_mask;
	wire [1:0] _readys_filter_T = ~readys_mask;
	wire [1:0] _readys_filter_T_1 = readys_valid & _readys_filter_T;
	wire [3:0] readys_filter = {_readys_filter_T_1, auto_out_1_d_valid, auto_out_0_d_valid};
	wire [3:0] _GEN_1 = {1'd0, readys_filter[3:1]};
	wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_1;
	wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0};
	wire [3:0] _GEN_2 = {1'd0, _readys_unready_T_1[3:1]};
	wire [3:0] readys_unready = _GEN_2 | _readys_unready_T_4;
	wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0];
	wire [1:0] readys_readys = ~_readys_readys_T_2;
	wire [1:0] _readys_mask_T = readys_readys & readys_valid;
	wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0};
	wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0];
	wire readys_0 = readys_readys[0];
	wire readys_1 = readys_readys[1];
	wire earlyWinner_0 = readys_0 & auto_out_0_d_valid;
	wire earlyWinner_1 = readys_1 & auto_out_1_d_valid;
	wire _prefixOR_T = earlyWinner_0 | earlyWinner_1;
	wire _T_10 = auto_out_0_d_valid | auto_out_1_d_valid;
	wire _T_11 = ~(auto_out_0_d_valid | auto_out_1_d_valid);
	reg state_0;
	wire muxStateEarly_0 = (idle ? earlyWinner_0 : state_0);
	reg state_1;
	wire muxStateEarly_1 = (idle ? earlyWinner_1 : state_1);
	wire _sink_ACancel_earlyValid_T_3 = (state_0 & auto_out_0_d_valid) | (state_1 & auto_out_1_d_valid);
	wire sink_ACancel_5_earlyValid = (idle ? _T_10 : _sink_ACancel_earlyValid_T_3);
	wire _beatsLeft_T_2 = auto_in_d_ready & sink_ACancel_5_earlyValid;
	wire allowed_0 = (idle ? readys_0 : state_0);
	wire allowed_1 = (idle ? readys_1 : state_1);
	wire [31:0] _T_27 = (muxStateEarly_0 ? auto_out_0_d_bits_data : 32'h00000000);
	wire [31:0] _T_28 = (muxStateEarly_1 ? auto_out_1_d_bits_data : 32'h00000000);
	wire [1:0] _T_39 = (muxStateEarly_0 ? auto_out_0_d_bits_size : 2'h0);
	wire [1:0] _T_40 = (muxStateEarly_1 ? 2'h2 : 2'h0);
	wire [2:0] _T_45 = (muxStateEarly_0 ? auto_out_0_d_bits_opcode : 3'h0);
	wire [2:0] _T_46 = (muxStateEarly_1 ? auto_out_1_d_bits_opcode : 3'h0);
	TLMonitor_36 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	assign auto_in_a_ready = (requestAIO_0_0 & auto_out_0_a_ready) | (requestAIO_0_1 & auto_out_1_a_ready);
	assign auto_in_d_valid = (idle ? _T_10 : _sink_ACancel_earlyValid_T_3);
	assign auto_in_d_bits_denied = muxStateEarly_0 & auto_out_0_d_bits_denied;
	assign auto_in_d_bits_data = _T_27 | _T_28;
	assign auto_in_d_bits_corrupt = muxStateEarly_0 & auto_out_0_d_bits_corrupt;
	assign auto_out_1_a_valid = auto_in_a_valid & requestAIO_0_1;
	assign auto_out_1_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_1_a_bits_address = auto_in_a_bits_address[6:0];
	assign auto_out_1_a_bits_data = auto_in_a_bits_data;
	assign auto_out_1_d_ready = auto_in_d_ready & allowed_1;
	assign auto_out_0_a_valid = auto_in_a_valid & requestAIO_0_0;
	assign auto_out_0_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_0_a_bits_address = auto_in_a_bits_address;
	assign auto_out_0_a_bits_data = auto_in_a_bits_data;
	assign auto_out_0_d_ready = auto_in_d_ready & allowed_0;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = (requestAIO_0_0 & auto_out_0_a_ready) | (requestAIO_0_1 & auto_out_1_a_ready);
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = (idle ? _T_10 : _sink_ACancel_earlyValid_T_3);
	assign monitor_io_in_d_bits_opcode = _T_45 | _T_46;
	assign monitor_io_in_d_bits_param = (muxStateEarly_0 ? auto_out_0_d_bits_param : 2'h0);
	assign monitor_io_in_d_bits_size = _T_39 | _T_40;
	assign monitor_io_in_d_bits_sink = muxStateEarly_0 & auto_out_0_d_bits_sink;
	assign monitor_io_in_d_bits_denied = muxStateEarly_0 & auto_out_0_d_bits_denied;
	assign monitor_io_in_d_bits_corrupt = muxStateEarly_0 & auto_out_0_d_bits_corrupt;
	always @(posedge clock) begin
		if (reset)
			beatsLeft <= 1'h0;
		else if (latch)
			beatsLeft <= 1'h0;
		else
			beatsLeft <= beatsLeft - _beatsLeft_T_2;
		if (reset)
			readys_mask <= 2'h3;
		else if (latch & |readys_valid)
			readys_mask <= _readys_mask_T_3;
		if (reset)
			state_0 <= 1'h0;
		else if (idle)
			state_0 <= earlyWinner_0;
		if (reset)
			state_1 <= 1'h0;
		else if (idle)
			state_1 <= earlyWinner_1;
	end
endmodule
module DMIToTL (
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_address,
	auto_out_a_bits_data,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt,
	io_dmi_req_ready,
	io_dmi_req_valid,
	io_dmi_req_bits_addr,
	io_dmi_req_bits_data,
	io_dmi_req_bits_op,
	io_dmi_resp_ready,
	io_dmi_resp_valid,
	io_dmi_resp_bits_data,
	io_dmi_resp_bits_resp
);
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [8:0] auto_out_a_bits_address;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input auto_out_d_bits_denied;
	input [31:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	output wire io_dmi_req_ready;
	input io_dmi_req_valid;
	input [6:0] io_dmi_req_bits_addr;
	input [31:0] io_dmi_req_bits_data;
	input [1:0] io_dmi_req_bits_op;
	input io_dmi_resp_ready;
	output wire io_dmi_resp_valid;
	output wire [31:0] io_dmi_resp_bits_data;
	output wire [1:0] io_dmi_resp_bits_resp;
	wire [8:0] addr = {io_dmi_req_bits_addr, 2'h0};
	wire [8:0] _GEN_3 = (io_dmi_req_bits_op == 2'h1 ? addr : 9'h048);
	wire [2:0] _GEN_7 = (io_dmi_req_bits_op == 2'h1 ? 3'h4 : 3'h0);
	wire _io_dmi_resp_bits_resp_T = auto_out_d_bits_corrupt | auto_out_d_bits_denied;
	assign auto_out_a_valid = io_dmi_req_valid;
	assign auto_out_a_bits_opcode = (io_dmi_req_bits_op == 2'h2 ? 3'h0 : _GEN_7);
	assign auto_out_a_bits_address = (io_dmi_req_bits_op == 2'h2 ? addr : _GEN_3);
	assign auto_out_a_bits_data = (io_dmi_req_bits_op == 2'h2 ? io_dmi_req_bits_data : 32'h00000000);
	assign auto_out_d_ready = io_dmi_resp_ready;
	assign io_dmi_req_ready = auto_out_a_ready;
	assign io_dmi_resp_valid = auto_out_d_valid;
	assign io_dmi_resp_bits_data = auto_out_d_bits_data;
	assign io_dmi_resp_bits_resp = {1'd0, _io_dmi_resp_bits_resp_T};
endmodule
module TLMonitor_37 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_address,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [6:0] io_in_a_bits_address;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire [6:0] _is_aligned_T = io_in_a_bits_address & 7'h03;
	wire is_aligned = _is_aligned_T == 7'h00;
	wire _T_15 = io_in_a_bits_opcode == 3'h6;
	wire [6:0] _T_20 = io_in_a_bits_address ^ 7'h40;
	wire [7:0] _T_21 = {1'b0, $signed(_T_20)};
	wire [7:0] _T_23 = $signed(_T_21) & -8'sh0c;
	wire _T_24 = $signed(_T_23) == 8'sh00;
	wire [6:0] _T_25 = io_in_a_bits_address ^ 7'h50;
	wire [7:0] _T_26 = {1'b0, $signed(_T_25)};
	wire [7:0] _T_28 = $signed(_T_26) & -8'sh08;
	wire _T_29 = $signed(_T_28) == 8'sh00;
	wire _T_30 = _T_24 | _T_29;
	wire _T_81 = io_in_a_bits_opcode == 3'h7;
	wire _T_151 = io_in_a_bits_opcode == 3'h4;
	wire _T_197 = io_in_a_bits_opcode == 3'h0;
	wire _T_237 = io_in_a_bits_opcode == 3'h1;
	wire _T_278 = io_in_a_bits_opcode == 3'h2;
	wire _T_314 = io_in_a_bits_opcode == 3'h3;
	wire _T_350 = io_in_a_bits_opcode == 3'h5;
	wire _T_390 = io_in_d_bits_opcode <= 3'h6;
	wire _T_394 = io_in_d_bits_opcode == 3'h6;
	wire _T_414 = io_in_d_bits_opcode == 3'h4;
	wire _T_442 = io_in_d_bits_opcode == 3'h5;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [6:0] address;
	wire _T_536 = io_in_a_valid & ~a_first;
	wire _T_537 = io_in_a_bits_opcode == opcode;
	wire _T_553 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	wire _T_560 = io_in_d_valid & ~d_first;
	wire _T_561 = io_in_d_bits_opcode == opcode_1;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [3:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_71 = {12'd0, inflight_opcodes};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_71 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [15:0] _GEN_73 = {12'd0, inflight_sizes};
	wire [15:0] _a_size_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_587 = io_in_a_valid & a_first_1;
	wire _T_590 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _a_opcodes_set_T_1 = {15'd0, a_opcodes_set_interm};
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? 3'h5 : 3'h0);
	wire [17:0] _a_sizes_set_T_1 = {15'd0, a_sizes_set_interm};
	wire _T_594 = ~inflight;
	wire [1:0] _GEN_16 = (a_first_done & a_first_1 ? 2'h1 : 2'h0);
	wire [18:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [17:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 18'h00000);
	wire _T_598 = io_in_d_valid & d_first_1;
	wire _T_600 = ~_T_394;
	wire _T_601 = (io_in_d_valid & d_first_1) & ~_T_394;
	wire [30:0] _d_opcodes_clr_T_5 = {15'd0, _a_opcode_lookup_T_5};
	wire [1:0] _GEN_22 = ((d_first_done & d_first_1) & _T_600 ? 2'h1 : 2'h0);
	wire [30:0] _GEN_23 = ((d_first_done & d_first_1) & _T_600 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire _T_613 = inflight | _T_587;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_618 = io_in_d_bits_opcode == _GEN_40;
	wire _T_619 = (io_in_d_bits_opcode == _GEN_32) | _T_618;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_630 = io_in_d_bits_opcode == _GEN_56;
	wire _T_631 = (io_in_d_bits_opcode == _GEN_48) | _T_630;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire _T_635 = 4'h2 == a_size_lookup;
	wire _T_645 = ((_T_598 & a_first_1) & io_in_a_valid) & _T_600;
	wire _T_647 = ~io_in_d_ready | io_in_a_ready;
	wire a_set = _GEN_16[0];
	wire d_clr = _GEN_22[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [3:0] a_sizes_set = _GEN_20[3:0];
	wire [3:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [3:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_656 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [3:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [15:0] _GEN_77 = {12'd0, inflight_sizes_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_77 & _a_opcode_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_682 = (io_in_d_valid & d_first_2) & _T_394;
	wire [30:0] _GEN_68 = ((d_first_done & d_first_2) & _T_394 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_700 = 4'h2 == c_size_lookup;
	wire [3:0] d_opcodes_clr_1 = _GEN_68[3:0];
	wire [3:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [3:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 4'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 4'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module TLDebugModuleOuter (
	clock,
	reset,
	auto_dmi_in_a_ready,
	auto_dmi_in_a_valid,
	auto_dmi_in_a_bits_opcode,
	auto_dmi_in_a_bits_address,
	auto_dmi_in_a_bits_data,
	auto_dmi_in_d_ready,
	auto_dmi_in_d_valid,
	auto_dmi_in_d_bits_opcode,
	auto_dmi_in_d_bits_data,
	auto_int_out_0,
	io_ctrl_dmactive,
	io_ctrl_dmactiveAck,
	io_innerCtrl_ready,
	io_innerCtrl_valid,
	io_innerCtrl_bits_resumereq,
	io_innerCtrl_bits_hartsel,
	io_innerCtrl_bits_ackhavereset,
	io_innerCtrl_bits_hrmask_0,
	io_hgDebugInt_0
);
	input clock;
	input reset;
	output wire auto_dmi_in_a_ready;
	input auto_dmi_in_a_valid;
	input [2:0] auto_dmi_in_a_bits_opcode;
	input [6:0] auto_dmi_in_a_bits_address;
	input [31:0] auto_dmi_in_a_bits_data;
	input auto_dmi_in_d_ready;
	output wire auto_dmi_in_d_valid;
	output wire [2:0] auto_dmi_in_d_bits_opcode;
	output wire [31:0] auto_dmi_in_d_bits_data;
	output wire auto_int_out_0;
	output wire io_ctrl_dmactive;
	input io_ctrl_dmactiveAck;
	input io_innerCtrl_ready;
	output wire io_innerCtrl_valid;
	output wire io_innerCtrl_bits_resumereq;
	output wire [9:0] io_innerCtrl_bits_hartsel;
	output wire io_innerCtrl_bits_ackhavereset;
	output wire io_innerCtrl_bits_hrmask_0;
	input io_hgDebugInt_0;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [6:0] monitor_io_in_a_bits_address;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	reg DMCONTROLReg_haltreq;
	reg DMCONTROLReg_ndmreset;
	reg DMCONTROLReg_dmactive;
	wire _T_1 = ~DMCONTROLReg_dmactive;
	wire in_bits_read = auto_dmi_in_a_bits_opcode == 3'h4;
	wire [2:0] in_bits_index = auto_dmi_in_a_bits_address[4:2];
	wire out_iindex = in_bits_index[1];
	wire [2:0] out_findex = in_bits_index & 3'h5;
	wire _out_T = out_findex == 3'h0;
	wire [1:0] _out_backSel_T = 2'h1 << out_iindex;
	wire out_backSel_0 = _out_backSel_T[0];
	wire out_woready_6 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_0) & (out_findex == 3'h0);
	wire DMCONTROLWrData_ndmreset = auto_dmi_in_a_bits_data[1];
	wire DMCONTROLWrData_haltreq = auto_dmi_in_a_bits_data[31];
	wire DMCONTROLWrData_dmactive = auto_dmi_in_a_bits_data[0];
	reg hrmaskReg_0;
	wire DMCONTROLWrData_clrresethaltreq = auto_dmi_in_a_bits_data[2];
	wire _T_11 = io_innerCtrl_bits_hartsel == 10'h000;
	wire DMCONTROLWrData_setresethaltreq = auto_dmi_in_a_bits_data[3];
	wire _GEN_23 = ((out_woready_6 & DMCONTROLWrData_setresethaltreq) & _T_11) | hrmaskReg_0;
	wire _GEN_24 = ((out_woready_6 & DMCONTROLWrData_clrresethaltreq) & _T_11 ? 1'h0 : _GEN_23);
	wire _T_18 = DMCONTROLReg_dmactive & io_ctrl_dmactiveAck;
	wire [4:0] out_prepend_7 = {3'h0, DMCONTROLReg_ndmreset, _T_18};
	wire [15:0] _out_T_96 = {11'd0, out_prepend_7};
	wire [17:0] out_prepend_9 = {2'h0, _out_T_96};
	wire [25:0] _out_T_114 = {8'd0, out_prepend_9};
	wire DMCONTROLWrData_ackhavereset = auto_dmi_in_a_bits_data[28];
	wire DMCONTROLWrData_resumereq = auto_dmi_in_a_bits_data[30];
	wire [31:0] out_prepend_15 = {DMCONTROLReg_haltreq, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, _out_T_114};
	wire _GEN_35 = (out_iindex ? _out_T : _out_T);
	wire [31:0] _GEN_37 = (out_iindex ? 32'h00111380 : out_prepend_15);
	reg debugIntRegs_0;
	reg innerCtrlValidReg;
	reg innerCtrlResumeReqReg;
	reg innerCtrlAckHaveResetReg;
	wire _innerCtrlValidReg_T = ~io_innerCtrl_ready;
	TLMonitor_37 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode)
	);
	assign auto_dmi_in_a_ready = auto_dmi_in_d_ready;
	assign auto_dmi_in_d_valid = auto_dmi_in_a_valid;
	assign auto_dmi_in_d_bits_opcode = {2'd0, in_bits_read};
	assign auto_dmi_in_d_bits_data = (_GEN_35 ? _GEN_37 : 32'h00000000);
	assign auto_int_out_0 = debugIntRegs_0 | io_hgDebugInt_0;
	assign io_ctrl_dmactive = DMCONTROLReg_dmactive;
	assign io_innerCtrl_valid = out_woready_6 | innerCtrlValidReg;
	assign io_innerCtrl_bits_resumereq = (out_woready_6 & DMCONTROLWrData_resumereq) | innerCtrlResumeReqReg;
	assign io_innerCtrl_bits_hartsel = 10'h000;
	assign io_innerCtrl_bits_ackhavereset = (out_woready_6 & DMCONTROLWrData_ackhavereset) | innerCtrlAckHaveResetReg;
	assign io_innerCtrl_bits_hrmask_0 = (_T_1 ? 1'h0 : _GEN_24);
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_dmi_in_d_ready;
	assign monitor_io_in_a_valid = auto_dmi_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_dmi_in_a_bits_opcode;
	assign monitor_io_in_a_bits_address = auto_dmi_in_a_bits_address;
	assign monitor_io_in_d_ready = auto_dmi_in_d_ready;
	assign monitor_io_in_d_valid = auto_dmi_in_a_valid;
	assign monitor_io_in_d_bits_opcode = {2'd0, in_bits_read};
	always @(posedge clock or posedge reset)
		if (reset)
			DMCONTROLReg_haltreq <= 1'h0;
		else if (~DMCONTROLReg_dmactive)
			DMCONTROLReg_haltreq <= 1'h0;
		else if (out_woready_6)
			DMCONTROLReg_haltreq <= DMCONTROLWrData_haltreq;
	always @(posedge clock or posedge reset)
		if (reset)
			DMCONTROLReg_ndmreset <= 1'h0;
		else if (~DMCONTROLReg_dmactive)
			DMCONTROLReg_ndmreset <= 1'h0;
		else if (out_woready_6)
			DMCONTROLReg_ndmreset <= DMCONTROLWrData_ndmreset;
	always @(posedge clock or posedge reset)
		if (reset)
			DMCONTROLReg_dmactive <= 1'h0;
		else if (out_woready_6)
			DMCONTROLReg_dmactive <= DMCONTROLWrData_dmactive;
		else if (~DMCONTROLReg_dmactive)
			DMCONTROLReg_dmactive <= 1'h0;
	always @(posedge clock or posedge reset)
		if (reset)
			hrmaskReg_0 <= 1'h0;
		else if (_T_1)
			hrmaskReg_0 <= 1'h0;
		else if ((out_woready_6 & DMCONTROLWrData_clrresethaltreq) & _T_11)
			hrmaskReg_0 <= 1'h0;
		else
			hrmaskReg_0 <= _GEN_23;
	always @(posedge clock or posedge reset)
		if (reset)
			debugIntRegs_0 <= 1'h0;
		else if (_T_1)
			debugIntRegs_0 <= 1'h0;
		else if (out_woready_6)
			debugIntRegs_0 <= DMCONTROLWrData_haltreq;
	always @(posedge clock or posedge reset)
		if (reset)
			innerCtrlValidReg <= 1'h0;
		else
			innerCtrlValidReg <= io_innerCtrl_valid & ~io_innerCtrl_ready;
	always @(posedge clock or posedge reset)
		if (reset)
			innerCtrlResumeReqReg <= 1'h0;
		else
			innerCtrlResumeReqReg <= io_innerCtrl_bits_resumereq & _innerCtrlValidReg_T;
	always @(posedge clock or posedge reset)
		if (reset)
			innerCtrlAckHaveResetReg <= 1'h0;
		else
			innerCtrlAckHaveResetReg <= io_innerCtrl_bits_ackhavereset & _innerCtrlValidReg_T;
endmodule
module IntSyncCrossingSource_4 (
	auto_in_0,
	auto_out_sync_0
);
	input auto_in_0;
	output wire auto_out_sync_0;
	assign auto_out_sync_0 = auto_in_0;
endmodule
module TLMonitor_38 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_address,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [8:0] io_in_a_bits_address;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [1:0] io_in_d_bits_size;
	input io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire [8:0] _is_aligned_T = io_in_a_bits_address & 9'h003;
	wire is_aligned = _is_aligned_T == 9'h000;
	wire [9:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_15 = io_in_a_bits_opcode == 3'h6;
	wire [9:0] _T_23 = $signed(_T_7) & -10'sh040;
	wire _T_24 = $signed(_T_23) == 10'sh000;
	wire [8:0] _T_25 = io_in_a_bits_address ^ 9'h044;
	wire [9:0] _T_26 = {1'b0, $signed(_T_25)};
	wire [9:0] _T_28 = $signed(_T_26) & -10'sh00c;
	wire _T_29 = $signed(_T_28) == 10'sh000;
	wire [8:0] _T_30 = io_in_a_bits_address ^ 9'h058;
	wire [9:0] _T_31 = {1'b0, $signed(_T_30)};
	wire [9:0] _T_33 = $signed(_T_31) & -10'sh008;
	wire _T_34 = $signed(_T_33) == 10'sh000;
	wire [8:0] _T_35 = io_in_a_bits_address ^ 9'h060;
	wire [9:0] _T_36 = {1'b0, $signed(_T_35)};
	wire [9:0] _T_38 = $signed(_T_36) & -10'sh020;
	wire _T_39 = $signed(_T_38) == 10'sh000;
	wire [8:0] _T_40 = io_in_a_bits_address ^ 9'h080;
	wire [9:0] _T_41 = {1'b0, $signed(_T_40)};
	wire [9:0] _T_43 = $signed(_T_41) & -10'sh080;
	wire _T_44 = $signed(_T_43) == 10'sh000;
	wire [8:0] _T_45 = io_in_a_bits_address ^ 9'h100;
	wire [9:0] _T_46 = {1'b0, $signed(_T_45)};
	wire [9:0] _T_48 = $signed(_T_46) & -10'sh100;
	wire _T_49 = $signed(_T_48) == 10'sh000;
	wire _T_54 = ((((_T_24 | _T_29) | _T_34) | _T_39) | _T_44) | _T_49;
	wire _T_129 = io_in_a_bits_opcode == 3'h7;
	wire _T_247 = io_in_a_bits_opcode == 3'h4;
	wire _T_317 = io_in_a_bits_opcode == 3'h0;
	wire _T_381 = io_in_a_bits_opcode == 3'h1;
	wire _T_446 = io_in_a_bits_opcode == 3'h2;
	wire _T_506 = io_in_a_bits_opcode == 3'h3;
	wire _T_566 = io_in_a_bits_opcode == 3'h5;
	wire _T_630 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_1 = ~io_in_d_bits_source;
	wire _T_634 = io_in_d_bits_opcode == 3'h6;
	wire _T_638 = io_in_d_bits_size >= 2'h2;
	wire _T_642 = io_in_d_bits_param == 2'h0;
	wire _T_646 = ~io_in_d_bits_corrupt;
	wire _T_650 = ~io_in_d_bits_denied;
	wire _T_654 = io_in_d_bits_opcode == 3'h4;
	wire _T_665 = io_in_d_bits_param <= 2'h2;
	wire _T_669 = io_in_d_bits_param != 2'h2;
	wire _T_682 = io_in_d_bits_opcode == 3'h5;
	wire _T_702 = _T_650 | io_in_d_bits_corrupt;
	wire _T_711 = io_in_d_bits_opcode == 3'h0;
	wire _T_728 = io_in_d_bits_opcode == 3'h1;
	wire _T_746 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [8:0] address;
	wire _T_776 = io_in_a_valid & ~a_first;
	wire _T_777 = io_in_a_bits_opcode == opcode;
	wire _T_793 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [1:0] size_1;
	reg source_1;
	reg sink;
	reg denied;
	wire _T_800 = io_in_d_valid & ~d_first;
	wire _T_801 = io_in_d_bits_opcode == opcode_1;
	wire _T_805 = io_in_d_bits_param == param_1;
	wire _T_809 = io_in_d_bits_size == size_1;
	wire _T_813 = io_in_d_bits_source == source_1;
	wire _T_817 = io_in_d_bits_sink == sink;
	wire _T_821 = io_in_d_bits_denied == denied;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [3:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [2:0] _GEN_71 = {io_in_d_bits_source, 2'h0};
	wire [3:0] _a_opcode_lookup_T = {1'd0, _GEN_71};
	wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_72 = {12'd0, _a_opcode_lookup_T_1};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_72 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [3:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [15:0] _GEN_75 = {12'd0, _a_size_lookup_T_1};
	wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_opcode_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_827 = io_in_a_valid & a_first_1;
	wire _T_830 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _a_opcodes_set_T_1 = {15'd0, a_opcodes_set_interm};
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? 3'h5 : 3'h0);
	wire [17:0] _a_sizes_set_T_1 = {15'd0, a_sizes_set_interm};
	wire _T_834 = ~inflight;
	wire [1:0] _GEN_16 = (a_first_done & a_first_1 ? 2'h1 : 2'h0);
	wire [18:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [17:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 18'h00000);
	wire _T_838 = io_in_d_valid & d_first_1;
	wire _T_840 = ~_T_634;
	wire _T_841 = (io_in_d_valid & d_first_1) & ~_T_634;
	wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source;
	wire [30:0] _GEN_1 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_opcodes_clr_T_5 = _GEN_1 << _a_opcode_lookup_T;
	wire [1:0] _GEN_22 = ((d_first_done & d_first_1) & _T_840 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_23 = ((d_first_done & d_first_1) & _T_840 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire same_cycle_resp = _T_827 & _source_ok_T_1;
	wire _T_853 = (inflight >> io_in_d_bits_source) | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_858 = io_in_d_bits_opcode == _GEN_40;
	wire _T_859 = (io_in_d_bits_opcode == _GEN_32) | _T_858;
	wire _T_863 = 2'h2 == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_870 = io_in_d_bits_opcode == _GEN_56;
	wire _T_871 = (io_in_d_bits_opcode == _GEN_48) | _T_870;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_79 = {2'd0, io_in_d_bits_size};
	wire _T_875 = _GEN_79 == a_size_lookup;
	wire _T_885 = (((_T_838 & a_first_1) & io_in_a_valid) & _source_ok_T_1) & _T_840;
	wire _T_887 = ~io_in_d_ready | io_in_a_ready;
	wire a_set = _GEN_16[0];
	wire d_clr = _GEN_22[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [3:0] a_sizes_set = _GEN_20[3:0];
	wire [3:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [3:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_896 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [3:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [3:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [15:0] _GEN_84 = {12'd0, _c_size_lookup_T_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_84 & _a_opcode_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_922 = (io_in_d_valid & d_first_2) & _T_634;
	wire [30:0] _GEN_68 = ((d_first_done & d_first_2) & _T_634 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire _T_930 = 1'h0 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_940 = _GEN_79 == c_size_lookup;
	wire [3:0] d_opcodes_clr_1 = _GEN_68[3:0];
	wire [3:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [3:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			param_1 <= io_in_d_bits_param;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (d_first_done & d_first)
			sink <= io_in_d_bits_sink;
		if (d_first_done & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 4'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 4'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module TLBusBypassBar (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_address,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_1_a_ready,
	auto_out_1_a_valid,
	auto_out_1_a_bits_opcode,
	auto_out_1_a_bits_address,
	auto_out_1_a_bits_data,
	auto_out_1_d_ready,
	auto_out_1_d_valid,
	auto_out_1_d_bits_opcode,
	auto_out_1_d_bits_param,
	auto_out_1_d_bits_size,
	auto_out_1_d_bits_source,
	auto_out_1_d_bits_sink,
	auto_out_1_d_bits_denied,
	auto_out_1_d_bits_data,
	auto_out_1_d_bits_corrupt,
	auto_out_0_a_ready,
	auto_out_0_a_valid,
	auto_out_0_a_bits_opcode,
	auto_out_0_a_bits_address,
	auto_out_0_d_ready,
	auto_out_0_d_valid,
	auto_out_0_d_bits_opcode,
	auto_out_0_d_bits_size,
	auto_out_0_d_bits_denied,
	auto_out_0_d_bits_corrupt,
	io_bypass
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [8:0] auto_in_a_bits_address;
	input [31:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [1:0] auto_in_d_bits_size;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_1_a_ready;
	output wire auto_out_1_a_valid;
	output wire [2:0] auto_out_1_a_bits_opcode;
	output wire [8:0] auto_out_1_a_bits_address;
	output wire [31:0] auto_out_1_a_bits_data;
	output wire auto_out_1_d_ready;
	input auto_out_1_d_valid;
	input [2:0] auto_out_1_d_bits_opcode;
	input [1:0] auto_out_1_d_bits_param;
	input [1:0] auto_out_1_d_bits_size;
	input auto_out_1_d_bits_source;
	input auto_out_1_d_bits_sink;
	input auto_out_1_d_bits_denied;
	input [31:0] auto_out_1_d_bits_data;
	input auto_out_1_d_bits_corrupt;
	input auto_out_0_a_ready;
	output wire auto_out_0_a_valid;
	output wire [2:0] auto_out_0_a_bits_opcode;
	output wire [127:0] auto_out_0_a_bits_address;
	output wire auto_out_0_d_ready;
	input auto_out_0_d_valid;
	input [2:0] auto_out_0_d_bits_opcode;
	input [1:0] auto_out_0_d_bits_size;
	input auto_out_0_d_bits_denied;
	input auto_out_0_d_bits_corrupt;
	input io_bypass;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [8:0] monitor_io_in_a_bits_address;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [1:0] monitor_io_in_d_bits_size;
	wire monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	reg in_reset;
	reg bypass_reg;
	wire bypass = (in_reset ? io_bypass : bypass_reg);
	reg [1:0] flight;
	reg stall_counter;
	wire stall_first = ~stall_counter;
	wire stall = (bypass != io_bypass) & stall_first;
	wire _bundleIn_0_a_ready_T = ~stall;
	wire _bundleIn_0_a_ready_T_1 = (bypass ? auto_out_0_a_ready : auto_out_1_a_ready);
	wire in_a_ready = ~stall & _bundleIn_0_a_ready_T_1;
	wire done = in_a_ready & auto_in_a_valid;
	reg counter;
	wire counter1 = counter - 1'h1;
	wire a_first = ~counter;
	wire in_d_valid = (bypass ? auto_out_0_d_valid : auto_out_1_d_valid);
	wire done_3 = auto_in_d_ready & in_d_valid;
	wire [2:0] in_d_bits_opcode = (bypass ? auto_out_0_d_bits_opcode : auto_out_1_d_bits_opcode);
	reg counter_3;
	wire counter1_3 = counter_3 - 1'h1;
	wire d_first = ~counter_3;
	wire d_request = in_d_bits_opcode[2] & ~in_d_bits_opcode[1];
	wire a_inc = done & a_first;
	wire d_inc = (done_3 & d_first) & d_request;
	wire [1:0] inc = {a_inc, d_inc};
	wire [1:0] dec = {1'h0, done_3};
	wire [1:0] _next_flight_T_2 = inc[0] + inc[1];
	wire [1:0] _next_flight_T_5 = flight + _next_flight_T_2;
	wire [1:0] _next_flight_T_8 = dec[0] + dec[1];
	wire [1:0] next_flight = _next_flight_T_5 - _next_flight_T_8;
	wire stall_counter1 = stall_counter - 1'h1;
	wire _bundleOut_0_a_valid_T_1 = _bundleIn_0_a_ready_T & auto_in_a_valid;
	wire _bundleOut_1_a_valid_T_2 = ~bypass;
	TLMonitor_38 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	assign auto_in_a_ready = ~stall & _bundleIn_0_a_ready_T_1;
	assign auto_in_d_valid = (bypass ? auto_out_0_d_valid : auto_out_1_d_valid);
	assign auto_in_d_bits_opcode = (bypass ? auto_out_0_d_bits_opcode : auto_out_1_d_bits_opcode);
	assign auto_in_d_bits_param = (bypass ? 2'h0 : auto_out_1_d_bits_param);
	assign auto_in_d_bits_size = (bypass ? auto_out_0_d_bits_size : auto_out_1_d_bits_size);
	assign auto_in_d_bits_sink = (bypass ? 1'h0 : auto_out_1_d_bits_sink);
	assign auto_in_d_bits_denied = (bypass ? auto_out_0_d_bits_denied : auto_out_1_d_bits_denied);
	assign auto_in_d_bits_data = (bypass ? 32'h00000000 : auto_out_1_d_bits_data);
	assign auto_in_d_bits_corrupt = (bypass ? auto_out_0_d_bits_corrupt : auto_out_1_d_bits_corrupt);
	assign auto_out_1_a_valid = _bundleOut_0_a_valid_T_1 & ~bypass;
	assign auto_out_1_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_1_a_bits_address = auto_in_a_bits_address;
	assign auto_out_1_a_bits_data = auto_in_a_bits_data;
	assign auto_out_1_d_ready = auto_in_d_ready & _bundleOut_1_a_valid_T_2;
	assign auto_out_0_a_valid = (_bundleIn_0_a_ready_T & auto_in_a_valid) & bypass;
	assign auto_out_0_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_0_a_bits_address = {119'd0, auto_in_a_bits_address};
	assign auto_out_0_d_ready = auto_in_d_ready & bypass;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = ~stall & _bundleIn_0_a_ready_T_1;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = (bypass ? auto_out_0_d_valid : auto_out_1_d_valid);
	assign monitor_io_in_d_bits_opcode = (bypass ? auto_out_0_d_bits_opcode : auto_out_1_d_bits_opcode);
	assign monitor_io_in_d_bits_param = (bypass ? 2'h0 : auto_out_1_d_bits_param);
	assign monitor_io_in_d_bits_size = (bypass ? auto_out_0_d_bits_size : auto_out_1_d_bits_size);
	assign monitor_io_in_d_bits_source = (bypass ? 1'h0 : auto_out_1_d_bits_source);
	assign monitor_io_in_d_bits_sink = (bypass ? 1'h0 : auto_out_1_d_bits_sink);
	assign monitor_io_in_d_bits_denied = (bypass ? auto_out_0_d_bits_denied : auto_out_1_d_bits_denied);
	assign monitor_io_in_d_bits_corrupt = (bypass ? auto_out_0_d_bits_corrupt : auto_out_1_d_bits_corrupt);
	always @(posedge clock) begin
		in_reset <= reset;
		if (in_reset | (next_flight == 2'h0))
			bypass_reg <= io_bypass;
		if (reset)
			flight <= 2'h0;
		else
			flight <= next_flight;
		if (reset)
			stall_counter <= 1'h0;
		else if (done)
			if (stall_first)
				stall_counter <= 1'h0;
			else
				stall_counter <= stall_counter1;
		if (reset)
			counter <= 1'h0;
		else if (done)
			if (a_first)
				counter <= 1'h0;
			else
				counter <= counter1;
		if (reset)
			counter_3 <= 1'h0;
		else if (done_3)
			if (d_first)
				counter_3 <= 1'h0;
			else
				counter_3 <= counter1_3;
	end
endmodule
module TLMonitor_39 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_address,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [127:0] io_in_a_bits_address;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_size;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire [127:0] _is_aligned_T = io_in_a_bits_address & 128'h00000000000000000000000000000003;
	wire is_aligned = _is_aligned_T == 128'h00000000000000000000000000000000;
	wire [128:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_15 = io_in_a_bits_opcode == 3'h6;
	wire [128:0] _T_26 = $signed(_T_7) & 129'sh100000000000000000000000000000000;
	wire _T_27 = $signed(_T_26) == 129'sh000000000000000000000000000000000;
	wire _T_72 = io_in_a_bits_opcode == 3'h7;
	wire _T_133 = io_in_a_bits_opcode == 3'h4;
	wire _T_173 = io_in_a_bits_opcode == 3'h0;
	wire _T_207 = io_in_a_bits_opcode == 3'h1;
	wire _T_242 = io_in_a_bits_opcode == 3'h2;
	wire _T_272 = io_in_a_bits_opcode == 3'h3;
	wire _T_302 = io_in_a_bits_opcode == 3'h5;
	wire _T_339 = io_in_d_bits_opcode <= 3'h6;
	wire _T_343 = io_in_d_bits_opcode == 3'h6;
	wire _T_347 = io_in_d_bits_size >= 2'h2;
	wire _T_355 = ~io_in_d_bits_corrupt;
	wire _T_359 = ~io_in_d_bits_denied;
	wire _T_363 = io_in_d_bits_opcode == 3'h4;
	wire _T_391 = io_in_d_bits_opcode == 3'h5;
	wire _T_411 = _T_359 | io_in_d_bits_corrupt;
	wire _T_420 = io_in_d_bits_opcode == 3'h0;
	wire _T_437 = io_in_d_bits_opcode == 3'h1;
	wire _T_455 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [127:0] address;
	wire _T_485 = io_in_a_valid & ~a_first;
	wire _T_486 = io_in_a_bits_opcode == opcode;
	wire _T_502 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] size_1;
	reg denied;
	wire _T_509 = io_in_d_valid & ~d_first;
	wire _T_510 = io_in_d_bits_opcode == opcode_1;
	wire _T_518 = io_in_d_bits_size == size_1;
	wire _T_530 = io_in_d_bits_denied == denied;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [3:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_71 = {12'd0, inflight_opcodes};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_71 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [15:0] _GEN_73 = {12'd0, inflight_sizes};
	wire [15:0] _a_size_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_536 = io_in_a_valid & a_first_1;
	wire _T_539 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _a_opcodes_set_T_1 = {15'd0, a_opcodes_set_interm};
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? 3'h5 : 3'h0);
	wire [17:0] _a_sizes_set_T_1 = {15'd0, a_sizes_set_interm};
	wire _T_543 = ~inflight;
	wire [1:0] _GEN_16 = (a_first_done & a_first_1 ? 2'h1 : 2'h0);
	wire [18:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [17:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 18'h00000);
	wire _T_547 = io_in_d_valid & d_first_1;
	wire _T_549 = ~_T_343;
	wire _T_550 = (io_in_d_valid & d_first_1) & ~_T_343;
	wire [30:0] _d_opcodes_clr_T_5 = {15'd0, _a_opcode_lookup_T_5};
	wire [1:0] _GEN_22 = ((d_first_done & d_first_1) & _T_549 ? 2'h1 : 2'h0);
	wire [30:0] _GEN_23 = ((d_first_done & d_first_1) & _T_549 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire _T_562 = inflight | _T_536;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_567 = io_in_d_bits_opcode == _GEN_40;
	wire _T_568 = (io_in_d_bits_opcode == _GEN_32) | _T_567;
	wire _T_572 = 2'h2 == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_579 = io_in_d_bits_opcode == _GEN_56;
	wire _T_580 = (io_in_d_bits_opcode == _GEN_48) | _T_579;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_75 = {2'd0, io_in_d_bits_size};
	wire _T_584 = _GEN_75 == a_size_lookup;
	wire _T_594 = ((_T_547 & a_first_1) & io_in_a_valid) & _T_549;
	wire _T_596 = ~io_in_d_ready | io_in_a_ready;
	wire a_set = _GEN_16[0];
	wire d_clr = _GEN_22[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [3:0] a_sizes_set = _GEN_20[3:0];
	wire [3:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [3:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_605 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [3:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [15:0] _GEN_78 = {12'd0, inflight_sizes_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_78 & _a_opcode_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_631 = (io_in_d_valid & d_first_2) & _T_343;
	wire [30:0] _GEN_68 = ((d_first_done & d_first_2) & _T_343 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_649 = _GEN_75 == c_size_lookup;
	wire [3:0] d_opcodes_clr_1 = _GEN_68[3:0];
	wire [3:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [3:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 4'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 4'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module TLError_1 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_address,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_denied,
	auto_in_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [127:0] auto_in_a_bits_address;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_size;
	output wire auto_in_d_bits_denied;
	output wire auto_in_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [127:0] monitor_io_in_a_bits_address;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_size;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	reg idle;
	reg beatsLeft;
	wire idle_1 = ~beatsLeft;
	wire da_valid = auto_in_a_valid & idle;
	wire [1:0] _readys_T = {da_valid, 1'h0};
	wire [2:0] _readys_T_1 = {_readys_T, 1'h0};
	wire [1:0] _readys_T_3 = _readys_T | _readys_T_1[1:0];
	wire [2:0] _readys_T_5 = {_readys_T_3, 1'h0};
	wire [1:0] _readys_T_7 = ~_readys_T_5[1:0];
	wire readys_1 = _readys_T_7[1];
	reg state_1;
	wire allowed_1 = (idle_1 ? readys_1 : state_1);
	wire out_1_ready = auto_in_d_ready & allowed_1;
	reg counter;
	wire [2:0] _GEN_4 = (3'h2 == auto_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_5 = (3'h3 == auto_in_a_bits_opcode ? 3'h1 : _GEN_4);
	wire [2:0] _GEN_6 = (3'h4 == auto_in_a_bits_opcode ? 3'h1 : _GEN_5);
	wire [2:0] _GEN_7 = (3'h5 == auto_in_a_bits_opcode ? 3'h2 : _GEN_6);
	wire [2:0] _GEN_8 = (3'h6 == auto_in_a_bits_opcode ? 3'h4 : _GEN_7);
	wire [2:0] da_bits_opcode = (3'h7 == auto_in_a_bits_opcode ? 3'h4 : _GEN_8);
	wire beats1_opdata = da_bits_opcode[0];
	wire done = out_1_ready & da_valid;
	wire counter1 = counter - 1'h1;
	wire da_first = ~counter;
	wire _T_3 = ~reset;
	wire _GEN_12 = (done & (da_bits_opcode == 3'h4) ? 1'h0 : idle);
	wire latch = idle_1 & auto_in_d_ready;
	wire earlyWinner_1 = readys_1 & da_valid;
	wire _T_22 = ~da_valid;
	wire muxStateEarly_1 = (idle_1 ? earlyWinner_1 : state_1);
	wire _sink_ACancel_earlyValid_T_2 = state_1 & da_valid;
	wire sink_ACancel_earlyValid = (idle_1 ? da_valid : _sink_ACancel_earlyValid_T_2);
	wire _beatsLeft_T_2 = auto_in_d_ready & sink_ACancel_earlyValid;
	TLMonitor_39 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	assign auto_in_a_ready = out_1_ready & idle;
	assign auto_in_d_valid = (idle_1 ? da_valid : _sink_ACancel_earlyValid_T_2);
	assign auto_in_d_bits_opcode = (muxStateEarly_1 ? da_bits_opcode : 3'h0);
	assign auto_in_d_bits_size = (muxStateEarly_1 ? 2'h2 : 2'h0);
	assign auto_in_d_bits_denied = (idle_1 ? earlyWinner_1 : state_1);
	assign auto_in_d_bits_corrupt = muxStateEarly_1 & beats1_opdata;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = out_1_ready & idle;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = (idle_1 ? da_valid : _sink_ACancel_earlyValid_T_2);
	assign monitor_io_in_d_bits_opcode = (muxStateEarly_1 ? da_bits_opcode : 3'h0);
	assign monitor_io_in_d_bits_size = (muxStateEarly_1 ? 2'h2 : 2'h0);
	assign monitor_io_in_d_bits_denied = (idle_1 ? earlyWinner_1 : state_1);
	assign monitor_io_in_d_bits_corrupt = muxStateEarly_1 & beats1_opdata;
	always @(posedge clock) begin
		idle <= reset | _GEN_12;
		if (reset)
			beatsLeft <= 1'h0;
		else if (latch)
			beatsLeft <= 1'h0;
		else
			beatsLeft <= beatsLeft - _beatsLeft_T_2;
		if (reset)
			state_1 <= 1'h0;
		else if (idle_1)
			state_1 <= earlyWinner_1;
		if (reset)
			counter <= 1'h0;
		else if (done)
			if (da_first)
				counter <= 1'h0;
			else
				counter <= counter1;
	end
endmodule
module TLBusBypass (
	clock,
	reset,
	auto_node_out_out_a_ready,
	auto_node_out_out_a_valid,
	auto_node_out_out_a_bits_opcode,
	auto_node_out_out_a_bits_address,
	auto_node_out_out_a_bits_data,
	auto_node_out_out_d_ready,
	auto_node_out_out_d_valid,
	auto_node_out_out_d_bits_opcode,
	auto_node_out_out_d_bits_param,
	auto_node_out_out_d_bits_size,
	auto_node_out_out_d_bits_source,
	auto_node_out_out_d_bits_sink,
	auto_node_out_out_d_bits_denied,
	auto_node_out_out_d_bits_data,
	auto_node_out_out_d_bits_corrupt,
	auto_node_in_in_a_ready,
	auto_node_in_in_a_valid,
	auto_node_in_in_a_bits_opcode,
	auto_node_in_in_a_bits_address,
	auto_node_in_in_a_bits_data,
	auto_node_in_in_d_ready,
	auto_node_in_in_d_valid,
	auto_node_in_in_d_bits_opcode,
	auto_node_in_in_d_bits_param,
	auto_node_in_in_d_bits_size,
	auto_node_in_in_d_bits_sink,
	auto_node_in_in_d_bits_denied,
	auto_node_in_in_d_bits_data,
	auto_node_in_in_d_bits_corrupt,
	io_bypass
);
	input clock;
	input reset;
	input auto_node_out_out_a_ready;
	output wire auto_node_out_out_a_valid;
	output wire [2:0] auto_node_out_out_a_bits_opcode;
	output wire [8:0] auto_node_out_out_a_bits_address;
	output wire [31:0] auto_node_out_out_a_bits_data;
	output wire auto_node_out_out_d_ready;
	input auto_node_out_out_d_valid;
	input [2:0] auto_node_out_out_d_bits_opcode;
	input [1:0] auto_node_out_out_d_bits_param;
	input [1:0] auto_node_out_out_d_bits_size;
	input auto_node_out_out_d_bits_source;
	input auto_node_out_out_d_bits_sink;
	input auto_node_out_out_d_bits_denied;
	input [31:0] auto_node_out_out_d_bits_data;
	input auto_node_out_out_d_bits_corrupt;
	output wire auto_node_in_in_a_ready;
	input auto_node_in_in_a_valid;
	input [2:0] auto_node_in_in_a_bits_opcode;
	input [8:0] auto_node_in_in_a_bits_address;
	input [31:0] auto_node_in_in_a_bits_data;
	input auto_node_in_in_d_ready;
	output wire auto_node_in_in_d_valid;
	output wire [2:0] auto_node_in_in_d_bits_opcode;
	output wire [1:0] auto_node_in_in_d_bits_param;
	output wire [1:0] auto_node_in_in_d_bits_size;
	output wire auto_node_in_in_d_bits_sink;
	output wire auto_node_in_in_d_bits_denied;
	output wire [31:0] auto_node_in_in_d_bits_data;
	output wire auto_node_in_in_d_bits_corrupt;
	input io_bypass;
	wire bar_clock;
	wire bar_reset;
	wire bar_auto_in_a_ready;
	wire bar_auto_in_a_valid;
	wire [2:0] bar_auto_in_a_bits_opcode;
	wire [8:0] bar_auto_in_a_bits_address;
	wire [31:0] bar_auto_in_a_bits_data;
	wire bar_auto_in_d_ready;
	wire bar_auto_in_d_valid;
	wire [2:0] bar_auto_in_d_bits_opcode;
	wire [1:0] bar_auto_in_d_bits_param;
	wire [1:0] bar_auto_in_d_bits_size;
	wire bar_auto_in_d_bits_sink;
	wire bar_auto_in_d_bits_denied;
	wire [31:0] bar_auto_in_d_bits_data;
	wire bar_auto_in_d_bits_corrupt;
	wire bar_auto_out_1_a_ready;
	wire bar_auto_out_1_a_valid;
	wire [2:0] bar_auto_out_1_a_bits_opcode;
	wire [8:0] bar_auto_out_1_a_bits_address;
	wire [31:0] bar_auto_out_1_a_bits_data;
	wire bar_auto_out_1_d_ready;
	wire bar_auto_out_1_d_valid;
	wire [2:0] bar_auto_out_1_d_bits_opcode;
	wire [1:0] bar_auto_out_1_d_bits_param;
	wire [1:0] bar_auto_out_1_d_bits_size;
	wire bar_auto_out_1_d_bits_source;
	wire bar_auto_out_1_d_bits_sink;
	wire bar_auto_out_1_d_bits_denied;
	wire [31:0] bar_auto_out_1_d_bits_data;
	wire bar_auto_out_1_d_bits_corrupt;
	wire bar_auto_out_0_a_ready;
	wire bar_auto_out_0_a_valid;
	wire [2:0] bar_auto_out_0_a_bits_opcode;
	wire [127:0] bar_auto_out_0_a_bits_address;
	wire bar_auto_out_0_d_ready;
	wire bar_auto_out_0_d_valid;
	wire [2:0] bar_auto_out_0_d_bits_opcode;
	wire [1:0] bar_auto_out_0_d_bits_size;
	wire bar_auto_out_0_d_bits_denied;
	wire bar_auto_out_0_d_bits_corrupt;
	wire bar_io_bypass;
	wire error_clock;
	wire error_reset;
	wire error_auto_in_a_ready;
	wire error_auto_in_a_valid;
	wire [2:0] error_auto_in_a_bits_opcode;
	wire [127:0] error_auto_in_a_bits_address;
	wire error_auto_in_d_ready;
	wire error_auto_in_d_valid;
	wire [2:0] error_auto_in_d_bits_opcode;
	wire [1:0] error_auto_in_d_bits_size;
	wire error_auto_in_d_bits_denied;
	wire error_auto_in_d_bits_corrupt;
	TLBusBypassBar bar(
		.clock(bar_clock),
		.reset(bar_reset),
		.auto_in_a_ready(bar_auto_in_a_ready),
		.auto_in_a_valid(bar_auto_in_a_valid),
		.auto_in_a_bits_opcode(bar_auto_in_a_bits_opcode),
		.auto_in_a_bits_address(bar_auto_in_a_bits_address),
		.auto_in_a_bits_data(bar_auto_in_a_bits_data),
		.auto_in_d_ready(bar_auto_in_d_ready),
		.auto_in_d_valid(bar_auto_in_d_valid),
		.auto_in_d_bits_opcode(bar_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(bar_auto_in_d_bits_param),
		.auto_in_d_bits_size(bar_auto_in_d_bits_size),
		.auto_in_d_bits_sink(bar_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(bar_auto_in_d_bits_denied),
		.auto_in_d_bits_data(bar_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(bar_auto_in_d_bits_corrupt),
		.auto_out_1_a_ready(bar_auto_out_1_a_ready),
		.auto_out_1_a_valid(bar_auto_out_1_a_valid),
		.auto_out_1_a_bits_opcode(bar_auto_out_1_a_bits_opcode),
		.auto_out_1_a_bits_address(bar_auto_out_1_a_bits_address),
		.auto_out_1_a_bits_data(bar_auto_out_1_a_bits_data),
		.auto_out_1_d_ready(bar_auto_out_1_d_ready),
		.auto_out_1_d_valid(bar_auto_out_1_d_valid),
		.auto_out_1_d_bits_opcode(bar_auto_out_1_d_bits_opcode),
		.auto_out_1_d_bits_param(bar_auto_out_1_d_bits_param),
		.auto_out_1_d_bits_size(bar_auto_out_1_d_bits_size),
		.auto_out_1_d_bits_source(bar_auto_out_1_d_bits_source),
		.auto_out_1_d_bits_sink(bar_auto_out_1_d_bits_sink),
		.auto_out_1_d_bits_denied(bar_auto_out_1_d_bits_denied),
		.auto_out_1_d_bits_data(bar_auto_out_1_d_bits_data),
		.auto_out_1_d_bits_corrupt(bar_auto_out_1_d_bits_corrupt),
		.auto_out_0_a_ready(bar_auto_out_0_a_ready),
		.auto_out_0_a_valid(bar_auto_out_0_a_valid),
		.auto_out_0_a_bits_opcode(bar_auto_out_0_a_bits_opcode),
		.auto_out_0_a_bits_address(bar_auto_out_0_a_bits_address),
		.auto_out_0_d_ready(bar_auto_out_0_d_ready),
		.auto_out_0_d_valid(bar_auto_out_0_d_valid),
		.auto_out_0_d_bits_opcode(bar_auto_out_0_d_bits_opcode),
		.auto_out_0_d_bits_size(bar_auto_out_0_d_bits_size),
		.auto_out_0_d_bits_denied(bar_auto_out_0_d_bits_denied),
		.auto_out_0_d_bits_corrupt(bar_auto_out_0_d_bits_corrupt),
		.io_bypass(bar_io_bypass)
	);
	TLError_1 error(
		.clock(error_clock),
		.reset(error_reset),
		.auto_in_a_ready(error_auto_in_a_ready),
		.auto_in_a_valid(error_auto_in_a_valid),
		.auto_in_a_bits_opcode(error_auto_in_a_bits_opcode),
		.auto_in_a_bits_address(error_auto_in_a_bits_address),
		.auto_in_d_ready(error_auto_in_d_ready),
		.auto_in_d_valid(error_auto_in_d_valid),
		.auto_in_d_bits_opcode(error_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(error_auto_in_d_bits_size),
		.auto_in_d_bits_denied(error_auto_in_d_bits_denied),
		.auto_in_d_bits_corrupt(error_auto_in_d_bits_corrupt)
	);
	assign auto_node_out_out_a_valid = bar_auto_out_1_a_valid;
	assign auto_node_out_out_a_bits_opcode = bar_auto_out_1_a_bits_opcode;
	assign auto_node_out_out_a_bits_address = bar_auto_out_1_a_bits_address;
	assign auto_node_out_out_a_bits_data = bar_auto_out_1_a_bits_data;
	assign auto_node_out_out_d_ready = bar_auto_out_1_d_ready;
	assign auto_node_in_in_a_ready = bar_auto_in_a_ready;
	assign auto_node_in_in_d_valid = bar_auto_in_d_valid;
	assign auto_node_in_in_d_bits_opcode = bar_auto_in_d_bits_opcode;
	assign auto_node_in_in_d_bits_param = bar_auto_in_d_bits_param;
	assign auto_node_in_in_d_bits_size = bar_auto_in_d_bits_size;
	assign auto_node_in_in_d_bits_sink = bar_auto_in_d_bits_sink;
	assign auto_node_in_in_d_bits_denied = bar_auto_in_d_bits_denied;
	assign auto_node_in_in_d_bits_data = bar_auto_in_d_bits_data;
	assign auto_node_in_in_d_bits_corrupt = bar_auto_in_d_bits_corrupt;
	assign bar_clock = clock;
	assign bar_reset = reset;
	assign bar_auto_in_a_valid = auto_node_in_in_a_valid;
	assign bar_auto_in_a_bits_opcode = auto_node_in_in_a_bits_opcode;
	assign bar_auto_in_a_bits_address = auto_node_in_in_a_bits_address;
	assign bar_auto_in_a_bits_data = auto_node_in_in_a_bits_data;
	assign bar_auto_in_d_ready = auto_node_in_in_d_ready;
	assign bar_auto_out_1_a_ready = auto_node_out_out_a_ready;
	assign bar_auto_out_1_d_valid = auto_node_out_out_d_valid;
	assign bar_auto_out_1_d_bits_opcode = auto_node_out_out_d_bits_opcode;
	assign bar_auto_out_1_d_bits_param = auto_node_out_out_d_bits_param;
	assign bar_auto_out_1_d_bits_size = auto_node_out_out_d_bits_size;
	assign bar_auto_out_1_d_bits_source = auto_node_out_out_d_bits_source;
	assign bar_auto_out_1_d_bits_sink = auto_node_out_out_d_bits_sink;
	assign bar_auto_out_1_d_bits_denied = auto_node_out_out_d_bits_denied;
	assign bar_auto_out_1_d_bits_data = auto_node_out_out_d_bits_data;
	assign bar_auto_out_1_d_bits_corrupt = auto_node_out_out_d_bits_corrupt;
	assign bar_auto_out_0_a_ready = error_auto_in_a_ready;
	assign bar_auto_out_0_d_valid = error_auto_in_d_valid;
	assign bar_auto_out_0_d_bits_opcode = error_auto_in_d_bits_opcode;
	assign bar_auto_out_0_d_bits_size = error_auto_in_d_bits_size;
	assign bar_auto_out_0_d_bits_denied = error_auto_in_d_bits_denied;
	assign bar_auto_out_0_d_bits_corrupt = error_auto_in_d_bits_corrupt;
	assign bar_io_bypass = io_bypass;
	assign error_clock = clock;
	assign error_reset = reset;
	assign error_auto_in_a_valid = bar_auto_out_0_a_valid;
	assign error_auto_in_a_bits_opcode = bar_auto_out_0_a_bits_opcode;
	assign error_auto_in_a_bits_address = bar_auto_out_0_a_bits_address;
	assign error_auto_in_d_ready = bar_auto_out_0_d_ready;
endmodule
module TLMonitor_40 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_address,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [8:0] io_in_a_bits_address;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [1:0] io_in_d_bits_size;
	input io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire [8:0] _is_aligned_T = io_in_a_bits_address & 9'h003;
	wire is_aligned = _is_aligned_T == 9'h000;
	wire [9:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_15 = io_in_a_bits_opcode == 3'h6;
	wire [9:0] _T_23 = $signed(_T_7) & -10'sh040;
	wire _T_24 = $signed(_T_23) == 10'sh000;
	wire [8:0] _T_25 = io_in_a_bits_address ^ 9'h044;
	wire [9:0] _T_26 = {1'b0, $signed(_T_25)};
	wire [9:0] _T_28 = $signed(_T_26) & -10'sh00c;
	wire _T_29 = $signed(_T_28) == 10'sh000;
	wire [8:0] _T_30 = io_in_a_bits_address ^ 9'h058;
	wire [9:0] _T_31 = {1'b0, $signed(_T_30)};
	wire [9:0] _T_33 = $signed(_T_31) & -10'sh008;
	wire _T_34 = $signed(_T_33) == 10'sh000;
	wire [8:0] _T_35 = io_in_a_bits_address ^ 9'h060;
	wire [9:0] _T_36 = {1'b0, $signed(_T_35)};
	wire [9:0] _T_38 = $signed(_T_36) & -10'sh020;
	wire _T_39 = $signed(_T_38) == 10'sh000;
	wire [8:0] _T_40 = io_in_a_bits_address ^ 9'h080;
	wire [9:0] _T_41 = {1'b0, $signed(_T_40)};
	wire [9:0] _T_43 = $signed(_T_41) & -10'sh080;
	wire _T_44 = $signed(_T_43) == 10'sh000;
	wire [8:0] _T_45 = io_in_a_bits_address ^ 9'h100;
	wire [9:0] _T_46 = {1'b0, $signed(_T_45)};
	wire [9:0] _T_48 = $signed(_T_46) & -10'sh100;
	wire _T_49 = $signed(_T_48) == 10'sh000;
	wire _T_54 = ((((_T_24 | _T_29) | _T_34) | _T_39) | _T_44) | _T_49;
	wire _T_129 = io_in_a_bits_opcode == 3'h7;
	wire _T_247 = io_in_a_bits_opcode == 3'h4;
	wire _T_317 = io_in_a_bits_opcode == 3'h0;
	wire _T_381 = io_in_a_bits_opcode == 3'h1;
	wire _T_446 = io_in_a_bits_opcode == 3'h2;
	wire _T_506 = io_in_a_bits_opcode == 3'h3;
	wire _T_566 = io_in_a_bits_opcode == 3'h5;
	wire _T_630 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_1 = ~io_in_d_bits_source;
	wire _T_634 = io_in_d_bits_opcode == 3'h6;
	wire _T_638 = io_in_d_bits_size >= 2'h2;
	wire _T_642 = io_in_d_bits_param == 2'h0;
	wire _T_646 = ~io_in_d_bits_corrupt;
	wire _T_650 = ~io_in_d_bits_denied;
	wire _T_654 = io_in_d_bits_opcode == 3'h4;
	wire _T_665 = io_in_d_bits_param <= 2'h2;
	wire _T_669 = io_in_d_bits_param != 2'h2;
	wire _T_682 = io_in_d_bits_opcode == 3'h5;
	wire _T_702 = _T_650 | io_in_d_bits_corrupt;
	wire _T_711 = io_in_d_bits_opcode == 3'h0;
	wire _T_728 = io_in_d_bits_opcode == 3'h1;
	wire _T_746 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [8:0] address;
	wire _T_776 = io_in_a_valid & ~a_first;
	wire _T_777 = io_in_a_bits_opcode == opcode;
	wire _T_793 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [1:0] size_1;
	reg source_1;
	reg sink;
	reg denied;
	wire _T_800 = io_in_d_valid & ~d_first;
	wire _T_801 = io_in_d_bits_opcode == opcode_1;
	wire _T_805 = io_in_d_bits_param == param_1;
	wire _T_809 = io_in_d_bits_size == size_1;
	wire _T_813 = io_in_d_bits_source == source_1;
	wire _T_817 = io_in_d_bits_sink == sink;
	wire _T_821 = io_in_d_bits_denied == denied;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [3:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [2:0] _GEN_71 = {io_in_d_bits_source, 2'h0};
	wire [3:0] _a_opcode_lookup_T = {1'd0, _GEN_71};
	wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_72 = {12'd0, _a_opcode_lookup_T_1};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_72 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [3:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [15:0] _GEN_75 = {12'd0, _a_size_lookup_T_1};
	wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_opcode_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_827 = io_in_a_valid & a_first_1;
	wire [1:0] _GEN_15 = (io_in_a_valid & a_first_1 ? 2'h1 : 2'h0);
	wire _T_830 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _a_opcodes_set_T_1 = {15'd0, a_opcodes_set_interm};
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? 3'h5 : 3'h0);
	wire [17:0] _a_sizes_set_T_1 = {15'd0, a_sizes_set_interm};
	wire _T_834 = ~inflight;
	wire [1:0] _GEN_16 = (a_first_done & a_first_1 ? 2'h1 : 2'h0);
	wire [18:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [17:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 18'h00000);
	wire _T_838 = io_in_d_valid & d_first_1;
	wire _T_840 = ~_T_634;
	wire _T_841 = (io_in_d_valid & d_first_1) & ~_T_634;
	wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source;
	wire [1:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_634 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_1 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_opcodes_clr_T_5 = _GEN_1 << _a_opcode_lookup_T;
	wire [1:0] _GEN_22 = ((d_first_done & d_first_1) & _T_840 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_23 = ((d_first_done & d_first_1) & _T_840 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire same_cycle_resp = _T_827 & _source_ok_T_1;
	wire _T_853 = (inflight >> io_in_d_bits_source) | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_858 = io_in_d_bits_opcode == _GEN_40;
	wire _T_859 = (io_in_d_bits_opcode == _GEN_32) | _T_858;
	wire _T_863 = 2'h2 == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_870 = io_in_d_bits_opcode == _GEN_56;
	wire _T_871 = (io_in_d_bits_opcode == _GEN_48) | _T_870;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_79 = {2'd0, io_in_d_bits_size};
	wire _T_875 = _GEN_79 == a_size_lookup;
	wire _T_885 = (((_T_838 & a_first_1) & io_in_a_valid) & _source_ok_T_1) & _T_840;
	wire _T_887 = ~io_in_d_ready | io_in_a_ready;
	wire a_set_wo_ready = _GEN_15[0];
	wire d_clr_wo_ready = _GEN_21[0];
	wire _T_894 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire a_set = _GEN_16[0];
	wire d_clr = _GEN_22[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [3:0] a_sizes_set = _GEN_20[3:0];
	wire [3:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [3:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_903 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [3:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [3:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [15:0] _GEN_84 = {12'd0, _c_size_lookup_T_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_84 & _a_opcode_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_929 = (io_in_d_valid & d_first_2) & _T_634;
	wire [30:0] _GEN_68 = ((d_first_done & d_first_2) & _T_634 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire _T_937 = 1'h0 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_947 = _GEN_79 == c_size_lookup;
	wire [3:0] d_opcodes_clr_1 = _GEN_68[3:0];
	wire [3:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [3:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			param_1 <= io_in_d_bits_param;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (d_first_done & d_first)
			sink <= io_in_d_bits_sink;
		if (d_first_done & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 4'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 4'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 (
	clock,
	reset,
	io_d,
	io_q
);
	input clock;
	input reset;
	input io_d;
	output wire io_q;
	reg sync_0;
	reg sync_1;
	reg sync_2;
	assign io_q = sync_0;
	always @(posedge clock or posedge reset)
		if (reset)
			sync_0 <= 1'h0;
		else
			sync_0 <= sync_1;
	always @(posedge clock or posedge reset)
		if (reset)
			sync_1 <= 1'h0;
		else
			sync_1 <= sync_2;
	always @(posedge clock or posedge reset)
		if (reset)
			sync_2 <= 1'h0;
		else
			sync_2 <= io_d;
endmodule
module AsyncResetSynchronizerShiftReg_w1_d3_i0 (
	clock,
	reset,
	io_d,
	io_q
);
	input clock;
	input reset;
	input io_d;
	output wire io_q;
	wire output_chain_clock;
	wire output_chain_reset;
	wire output_chain_io_d;
	wire output_chain_io_q;
	AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain(
		.clock(output_chain_clock),
		.reset(output_chain_reset),
		.io_d(output_chain_io_d),
		.io_q(output_chain_io_q)
	);
	assign io_q = output_chain_io_q;
	assign output_chain_clock = clock;
	assign output_chain_reset = reset;
	assign output_chain_io_d = io_d;
endmodule
module AsyncResetSynchronizerShiftReg_w1_d3_i0_1 (
	clock,
	reset,
	io_d,
	io_q
);
	input clock;
	input reset;
	input io_d;
	output wire io_q;
	wire output_chain_clock;
	wire output_chain_reset;
	wire output_chain_io_d;
	wire output_chain_io_q;
	AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain(
		.clock(output_chain_clock),
		.reset(output_chain_reset),
		.io_d(output_chain_io_d),
		.io_q(output_chain_io_q)
	);
	assign io_q = output_chain_io_q;
	assign output_chain_clock = clock;
	assign output_chain_reset = reset;
	assign output_chain_io_d = io_d;
endmodule
module AsyncValidSync (
	io_in,
	io_out,
	clock,
	reset
);
	input io_in;
	output wire io_out;
	input clock;
	input reset;
	wire io_out_source_valid_0_clock;
	wire io_out_source_valid_0_reset;
	wire io_out_source_valid_0_io_d;
	wire io_out_source_valid_0_io_q;
	AsyncResetSynchronizerShiftReg_w1_d3_i0_1 io_out_source_valid_0(
		.clock(io_out_source_valid_0_clock),
		.reset(io_out_source_valid_0_reset),
		.io_d(io_out_source_valid_0_io_d),
		.io_q(io_out_source_valid_0_io_q)
	);
	assign io_out = io_out_source_valid_0_io_q;
	assign io_out_source_valid_0_clock = clock;
	assign io_out_source_valid_0_reset = reset;
	assign io_out_source_valid_0_io_d = io_in;
endmodule
module AsyncQueueSource (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_address,
	io_enq_bits_data,
	io_async_mem_0_opcode,
	io_async_mem_0_address,
	io_async_mem_0_data,
	io_async_ridx,
	io_async_widx,
	io_async_safe_ridx_valid,
	io_async_safe_widx_valid,
	io_async_safe_source_reset_n,
	io_async_safe_sink_reset_n
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [8:0] io_enq_bits_address;
	input [31:0] io_enq_bits_data;
	output wire [2:0] io_async_mem_0_opcode;
	output wire [8:0] io_async_mem_0_address;
	output wire [31:0] io_async_mem_0_data;
	input io_async_ridx;
	output wire io_async_widx;
	input io_async_safe_ridx_valid;
	output wire io_async_safe_widx_valid;
	output wire io_async_safe_source_reset_n;
	input io_async_safe_sink_reset_n;
	wire ridx_ridx_gray_clock;
	wire ridx_ridx_gray_reset;
	wire ridx_ridx_gray_io_d;
	wire ridx_ridx_gray_io_q;
	wire source_valid_0_io_in;
	wire source_valid_0_io_out;
	wire source_valid_0_clock;
	wire source_valid_0_reset;
	wire source_valid_1_io_in;
	wire source_valid_1_io_out;
	wire source_valid_1_clock;
	wire source_valid_1_reset;
	wire sink_extend_io_in;
	wire sink_extend_io_out;
	wire sink_extend_clock;
	wire sink_extend_reset;
	wire sink_valid_io_in;
	wire sink_valid_io_out;
	wire sink_valid_clock;
	wire sink_valid_reset;
	reg [2:0] mem_0_opcode;
	reg [8:0] mem_0_address;
	reg [31:0] mem_0_data;
	wire _widx_T_1 = io_enq_ready & io_enq_valid;
	wire sink_ready = sink_valid_io_out;
	wire _widx_T_2 = ~sink_ready;
	reg widx_widx_bin;
	wire widx_incremented = (_widx_T_2 ? 1'h0 : widx_widx_bin + _widx_T_1);
	wire ridx = ridx_ridx_gray_io_q;
	reg ready_reg;
	reg widx_gray;
	AsyncResetSynchronizerShiftReg_w1_d3_i0 ridx_ridx_gray(
		.clock(ridx_ridx_gray_clock),
		.reset(ridx_ridx_gray_reset),
		.io_d(ridx_ridx_gray_io_d),
		.io_q(ridx_ridx_gray_io_q)
	);
	AsyncValidSync source_valid_0(
		.io_in(source_valid_0_io_in),
		.io_out(source_valid_0_io_out),
		.clock(source_valid_0_clock),
		.reset(source_valid_0_reset)
	);
	AsyncValidSync source_valid_1(
		.io_in(source_valid_1_io_in),
		.io_out(source_valid_1_io_out),
		.clock(source_valid_1_clock),
		.reset(source_valid_1_reset)
	);
	AsyncValidSync sink_extend(
		.io_in(sink_extend_io_in),
		.io_out(sink_extend_io_out),
		.clock(sink_extend_clock),
		.reset(sink_extend_reset)
	);
	AsyncValidSync sink_valid(
		.io_in(sink_valid_io_in),
		.io_out(sink_valid_io_out),
		.clock(sink_valid_clock),
		.reset(sink_valid_reset)
	);
	assign io_enq_ready = ready_reg & sink_ready;
	assign io_async_mem_0_opcode = mem_0_opcode;
	assign io_async_mem_0_address = mem_0_address;
	assign io_async_mem_0_data = mem_0_data;
	assign io_async_widx = widx_gray;
	assign io_async_safe_widx_valid = source_valid_1_io_out;
	assign io_async_safe_source_reset_n = ~reset;
	assign ridx_ridx_gray_clock = clock;
	assign ridx_ridx_gray_reset = reset;
	assign ridx_ridx_gray_io_d = io_async_ridx;
	assign source_valid_0_io_in = 1'h1;
	assign source_valid_0_clock = clock;
	assign source_valid_0_reset = reset | ~io_async_safe_sink_reset_n;
	assign source_valid_1_io_in = source_valid_0_io_out;
	assign source_valid_1_clock = clock;
	assign source_valid_1_reset = reset | ~io_async_safe_sink_reset_n;
	assign sink_extend_io_in = io_async_safe_ridx_valid;
	assign sink_extend_clock = clock;
	assign sink_extend_reset = reset | ~io_async_safe_sink_reset_n;
	assign sink_valid_io_in = sink_extend_io_out;
	assign sink_valid_clock = clock;
	assign sink_valid_reset = reset;
	always @(posedge clock) begin
		if (_widx_T_1)
			mem_0_opcode <= io_enq_bits_opcode;
		if (_widx_T_1)
			mem_0_address <= io_enq_bits_address;
		if (_widx_T_1)
			mem_0_data <= io_enq_bits_data;
	end
	always @(posedge clock or posedge reset)
		if (reset)
			widx_widx_bin <= 1'h0;
		else if (_widx_T_2)
			widx_widx_bin <= 1'h0;
		else
			widx_widx_bin <= widx_widx_bin + _widx_T_1;
	always @(posedge clock or posedge reset)
		if (reset)
			ready_reg <= 1'h0;
		else
			ready_reg <= sink_ready & (widx_incremented != (ridx ^ 1'h1));
	always @(posedge clock or posedge reset)
		if (reset)
			widx_gray <= 1'h0;
		else if (_widx_T_2)
			widx_gray <= 1'h0;
		else
			widx_gray <= widx_widx_bin + _widx_T_1;
endmodule
module ClockCrossingReg_w43 (
	clock,
	io_d,
	io_q,
	io_en
);
	input clock;
	input [42:0] io_d;
	output wire [42:0] io_q;
	input io_en;
	reg [42:0] cdc_reg;
	assign io_q = cdc_reg;
	always @(posedge clock)
		if (io_en)
			cdc_reg <= io_d;
endmodule
module AsyncQueueSink (
	clock,
	reset,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_sink,
	io_deq_bits_denied,
	io_deq_bits_data,
	io_deq_bits_corrupt,
	io_async_mem_0_opcode,
	io_async_mem_0_size,
	io_async_mem_0_source,
	io_async_mem_0_data,
	io_async_ridx,
	io_async_widx,
	io_async_safe_ridx_valid,
	io_async_safe_widx_valid,
	io_async_safe_source_reset_n,
	io_async_safe_sink_reset_n
);
	input clock;
	input reset;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [1:0] io_deq_bits_param;
	output wire [1:0] io_deq_bits_size;
	output wire io_deq_bits_source;
	output wire io_deq_bits_sink;
	output wire io_deq_bits_denied;
	output wire [31:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	input [2:0] io_async_mem_0_opcode;
	input [1:0] io_async_mem_0_size;
	input io_async_mem_0_source;
	input [31:0] io_async_mem_0_data;
	output wire io_async_ridx;
	input io_async_widx;
	output wire io_async_safe_ridx_valid;
	input io_async_safe_widx_valid;
	input io_async_safe_source_reset_n;
	output wire io_async_safe_sink_reset_n;
	wire widx_widx_gray_clock;
	wire widx_widx_gray_reset;
	wire widx_widx_gray_io_d;
	wire widx_widx_gray_io_q;
	wire io_deq_bits_deq_bits_reg_clock;
	wire [42:0] io_deq_bits_deq_bits_reg_io_d;
	wire [42:0] io_deq_bits_deq_bits_reg_io_q;
	wire io_deq_bits_deq_bits_reg_io_en;
	wire sink_valid_0_io_in;
	wire sink_valid_0_io_out;
	wire sink_valid_0_clock;
	wire sink_valid_0_reset;
	wire sink_valid_1_io_in;
	wire sink_valid_1_io_out;
	wire sink_valid_1_clock;
	wire sink_valid_1_reset;
	wire source_extend_io_in;
	wire source_extend_io_out;
	wire source_extend_clock;
	wire source_extend_reset;
	wire source_valid_io_in;
	wire source_valid_io_out;
	wire source_valid_clock;
	wire source_valid_reset;
	wire _ridx_T_1 = io_deq_ready & io_deq_valid;
	wire source_ready = source_valid_io_out;
	wire _ridx_T_2 = ~source_ready;
	reg ridx_ridx_bin;
	wire ridx_incremented = (_ridx_T_2 ? 1'h0 : ridx_ridx_bin + _ridx_T_1);
	wire widx = widx_widx_gray_io_q;
	wire [34:0] io_deq_bits_deq_bits_reg_io_d_lo = {2'h0, io_async_mem_0_data, 1'h0};
	wire [7:0] io_deq_bits_deq_bits_reg_io_d_hi = {io_async_mem_0_opcode, 2'h0, io_async_mem_0_size, io_async_mem_0_source};
	wire [42:0] _io_deq_bits_WIRE_1 = io_deq_bits_deq_bits_reg_io_q;
	reg valid_reg;
	reg ridx_gray;
	AsyncResetSynchronizerShiftReg_w1_d3_i0 widx_widx_gray(
		.clock(widx_widx_gray_clock),
		.reset(widx_widx_gray_reset),
		.io_d(widx_widx_gray_io_d),
		.io_q(widx_widx_gray_io_q)
	);
	ClockCrossingReg_w43 io_deq_bits_deq_bits_reg(
		.clock(io_deq_bits_deq_bits_reg_clock),
		.io_d(io_deq_bits_deq_bits_reg_io_d),
		.io_q(io_deq_bits_deq_bits_reg_io_q),
		.io_en(io_deq_bits_deq_bits_reg_io_en)
	);
	AsyncValidSync sink_valid_0(
		.io_in(sink_valid_0_io_in),
		.io_out(sink_valid_0_io_out),
		.clock(sink_valid_0_clock),
		.reset(sink_valid_0_reset)
	);
	AsyncValidSync sink_valid_1(
		.io_in(sink_valid_1_io_in),
		.io_out(sink_valid_1_io_out),
		.clock(sink_valid_1_clock),
		.reset(sink_valid_1_reset)
	);
	AsyncValidSync source_extend(
		.io_in(source_extend_io_in),
		.io_out(source_extend_io_out),
		.clock(source_extend_clock),
		.reset(source_extend_reset)
	);
	AsyncValidSync source_valid(
		.io_in(source_valid_io_in),
		.io_out(source_valid_io_out),
		.clock(source_valid_clock),
		.reset(source_valid_reset)
	);
	assign io_deq_valid = valid_reg & source_ready;
	assign io_deq_bits_opcode = _io_deq_bits_WIRE_1[42:40];
	assign io_deq_bits_param = _io_deq_bits_WIRE_1[39:38];
	assign io_deq_bits_size = _io_deq_bits_WIRE_1[37:36];
	assign io_deq_bits_source = _io_deq_bits_WIRE_1[35];
	assign io_deq_bits_sink = _io_deq_bits_WIRE_1[34];
	assign io_deq_bits_denied = _io_deq_bits_WIRE_1[33];
	assign io_deq_bits_data = _io_deq_bits_WIRE_1[32:1];
	assign io_deq_bits_corrupt = _io_deq_bits_WIRE_1[0];
	assign io_async_ridx = ridx_gray;
	assign io_async_safe_ridx_valid = sink_valid_1_io_out;
	assign io_async_safe_sink_reset_n = ~reset;
	assign widx_widx_gray_clock = clock;
	assign widx_widx_gray_reset = reset;
	assign widx_widx_gray_io_d = io_async_widx;
	assign io_deq_bits_deq_bits_reg_clock = clock;
	assign io_deq_bits_deq_bits_reg_io_d = {io_deq_bits_deq_bits_reg_io_d_hi, io_deq_bits_deq_bits_reg_io_d_lo};
	assign io_deq_bits_deq_bits_reg_io_en = source_ready & (ridx_incremented != widx);
	assign sink_valid_0_io_in = 1'h1;
	assign sink_valid_0_clock = clock;
	assign sink_valid_0_reset = reset | ~io_async_safe_source_reset_n;
	assign sink_valid_1_io_in = sink_valid_0_io_out;
	assign sink_valid_1_clock = clock;
	assign sink_valid_1_reset = reset | ~io_async_safe_source_reset_n;
	assign source_extend_io_in = io_async_safe_widx_valid;
	assign source_extend_clock = clock;
	assign source_extend_reset = reset | ~io_async_safe_source_reset_n;
	assign source_valid_io_in = source_extend_io_out;
	assign source_valid_clock = clock;
	assign source_valid_reset = reset;
	always @(posedge clock or posedge reset)
		if (reset)
			ridx_ridx_bin <= 1'h0;
		else if (_ridx_T_2)
			ridx_ridx_bin <= 1'h0;
		else
			ridx_ridx_bin <= ridx_ridx_bin + _ridx_T_1;
	always @(posedge clock or posedge reset)
		if (reset)
			valid_reg <= 1'h0;
		else
			valid_reg <= source_ready & (ridx_incremented != widx);
	always @(posedge clock or posedge reset)
		if (reset)
			ridx_gray <= 1'h0;
		else if (_ridx_T_2)
			ridx_gray <= 1'h0;
		else
			ridx_gray <= ridx_ridx_bin + _ridx_T_1;
endmodule
module TLAsyncCrossingSource (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_address,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_mem_0_opcode,
	auto_out_a_mem_0_address,
	auto_out_a_mem_0_data,
	auto_out_a_ridx,
	auto_out_a_widx,
	auto_out_a_safe_ridx_valid,
	auto_out_a_safe_widx_valid,
	auto_out_a_safe_source_reset_n,
	auto_out_a_safe_sink_reset_n,
	auto_out_d_mem_0_opcode,
	auto_out_d_mem_0_size,
	auto_out_d_mem_0_source,
	auto_out_d_mem_0_data,
	auto_out_d_ridx,
	auto_out_d_widx,
	auto_out_d_safe_ridx_valid,
	auto_out_d_safe_widx_valid,
	auto_out_d_safe_source_reset_n,
	auto_out_d_safe_sink_reset_n
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [8:0] auto_in_a_bits_address;
	input [31:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [1:0] auto_in_d_bits_size;
	output wire auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [31:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	output wire [2:0] auto_out_a_mem_0_opcode;
	output wire [8:0] auto_out_a_mem_0_address;
	output wire [31:0] auto_out_a_mem_0_data;
	input auto_out_a_ridx;
	output wire auto_out_a_widx;
	input auto_out_a_safe_ridx_valid;
	output wire auto_out_a_safe_widx_valid;
	output wire auto_out_a_safe_source_reset_n;
	input auto_out_a_safe_sink_reset_n;
	input [2:0] auto_out_d_mem_0_opcode;
	input [1:0] auto_out_d_mem_0_size;
	input auto_out_d_mem_0_source;
	input [31:0] auto_out_d_mem_0_data;
	output wire auto_out_d_ridx;
	input auto_out_d_widx;
	output wire auto_out_d_safe_ridx_valid;
	input auto_out_d_safe_widx_valid;
	input auto_out_d_safe_source_reset_n;
	output wire auto_out_d_safe_sink_reset_n;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [8:0] monitor_io_in_a_bits_address;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [1:0] monitor_io_in_d_bits_size;
	wire monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire bundleOut_0_a_source_clock;
	wire bundleOut_0_a_source_reset;
	wire bundleOut_0_a_source_io_enq_ready;
	wire bundleOut_0_a_source_io_enq_valid;
	wire [2:0] bundleOut_0_a_source_io_enq_bits_opcode;
	wire [8:0] bundleOut_0_a_source_io_enq_bits_address;
	wire [31:0] bundleOut_0_a_source_io_enq_bits_data;
	wire [2:0] bundleOut_0_a_source_io_async_mem_0_opcode;
	wire [8:0] bundleOut_0_a_source_io_async_mem_0_address;
	wire [31:0] bundleOut_0_a_source_io_async_mem_0_data;
	wire bundleOut_0_a_source_io_async_ridx;
	wire bundleOut_0_a_source_io_async_widx;
	wire bundleOut_0_a_source_io_async_safe_ridx_valid;
	wire bundleOut_0_a_source_io_async_safe_widx_valid;
	wire bundleOut_0_a_source_io_async_safe_source_reset_n;
	wire bundleOut_0_a_source_io_async_safe_sink_reset_n;
	wire bundleIn_0_d_sink_clock;
	wire bundleIn_0_d_sink_reset;
	wire bundleIn_0_d_sink_io_deq_ready;
	wire bundleIn_0_d_sink_io_deq_valid;
	wire [2:0] bundleIn_0_d_sink_io_deq_bits_opcode;
	wire [1:0] bundleIn_0_d_sink_io_deq_bits_param;
	wire [1:0] bundleIn_0_d_sink_io_deq_bits_size;
	wire bundleIn_0_d_sink_io_deq_bits_source;
	wire bundleIn_0_d_sink_io_deq_bits_sink;
	wire bundleIn_0_d_sink_io_deq_bits_denied;
	wire [31:0] bundleIn_0_d_sink_io_deq_bits_data;
	wire bundleIn_0_d_sink_io_deq_bits_corrupt;
	wire [2:0] bundleIn_0_d_sink_io_async_mem_0_opcode;
	wire [1:0] bundleIn_0_d_sink_io_async_mem_0_size;
	wire bundleIn_0_d_sink_io_async_mem_0_source;
	wire [31:0] bundleIn_0_d_sink_io_async_mem_0_data;
	wire bundleIn_0_d_sink_io_async_ridx;
	wire bundleIn_0_d_sink_io_async_widx;
	wire bundleIn_0_d_sink_io_async_safe_ridx_valid;
	wire bundleIn_0_d_sink_io_async_safe_widx_valid;
	wire bundleIn_0_d_sink_io_async_safe_source_reset_n;
	wire bundleIn_0_d_sink_io_async_safe_sink_reset_n;
	TLMonitor_40 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	AsyncQueueSource bundleOut_0_a_source(
		.clock(bundleOut_0_a_source_clock),
		.reset(bundleOut_0_a_source_reset),
		.io_enq_ready(bundleOut_0_a_source_io_enq_ready),
		.io_enq_valid(bundleOut_0_a_source_io_enq_valid),
		.io_enq_bits_opcode(bundleOut_0_a_source_io_enq_bits_opcode),
		.io_enq_bits_address(bundleOut_0_a_source_io_enq_bits_address),
		.io_enq_bits_data(bundleOut_0_a_source_io_enq_bits_data),
		.io_async_mem_0_opcode(bundleOut_0_a_source_io_async_mem_0_opcode),
		.io_async_mem_0_address(bundleOut_0_a_source_io_async_mem_0_address),
		.io_async_mem_0_data(bundleOut_0_a_source_io_async_mem_0_data),
		.io_async_ridx(bundleOut_0_a_source_io_async_ridx),
		.io_async_widx(bundleOut_0_a_source_io_async_widx),
		.io_async_safe_ridx_valid(bundleOut_0_a_source_io_async_safe_ridx_valid),
		.io_async_safe_widx_valid(bundleOut_0_a_source_io_async_safe_widx_valid),
		.io_async_safe_source_reset_n(bundleOut_0_a_source_io_async_safe_source_reset_n),
		.io_async_safe_sink_reset_n(bundleOut_0_a_source_io_async_safe_sink_reset_n)
	);
	AsyncQueueSink bundleIn_0_d_sink(
		.clock(bundleIn_0_d_sink_clock),
		.reset(bundleIn_0_d_sink_reset),
		.io_deq_ready(bundleIn_0_d_sink_io_deq_ready),
		.io_deq_valid(bundleIn_0_d_sink_io_deq_valid),
		.io_deq_bits_opcode(bundleIn_0_d_sink_io_deq_bits_opcode),
		.io_deq_bits_param(bundleIn_0_d_sink_io_deq_bits_param),
		.io_deq_bits_size(bundleIn_0_d_sink_io_deq_bits_size),
		.io_deq_bits_source(bundleIn_0_d_sink_io_deq_bits_source),
		.io_deq_bits_sink(bundleIn_0_d_sink_io_deq_bits_sink),
		.io_deq_bits_denied(bundleIn_0_d_sink_io_deq_bits_denied),
		.io_deq_bits_data(bundleIn_0_d_sink_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleIn_0_d_sink_io_deq_bits_corrupt),
		.io_async_mem_0_opcode(bundleIn_0_d_sink_io_async_mem_0_opcode),
		.io_async_mem_0_size(bundleIn_0_d_sink_io_async_mem_0_size),
		.io_async_mem_0_source(bundleIn_0_d_sink_io_async_mem_0_source),
		.io_async_mem_0_data(bundleIn_0_d_sink_io_async_mem_0_data),
		.io_async_ridx(bundleIn_0_d_sink_io_async_ridx),
		.io_async_widx(bundleIn_0_d_sink_io_async_widx),
		.io_async_safe_ridx_valid(bundleIn_0_d_sink_io_async_safe_ridx_valid),
		.io_async_safe_widx_valid(bundleIn_0_d_sink_io_async_safe_widx_valid),
		.io_async_safe_source_reset_n(bundleIn_0_d_sink_io_async_safe_source_reset_n),
		.io_async_safe_sink_reset_n(bundleIn_0_d_sink_io_async_safe_sink_reset_n)
	);
	assign auto_in_a_ready = bundleOut_0_a_source_io_enq_ready;
	assign auto_in_d_valid = bundleIn_0_d_sink_io_deq_valid;
	assign auto_in_d_bits_opcode = bundleIn_0_d_sink_io_deq_bits_opcode;
	assign auto_in_d_bits_param = bundleIn_0_d_sink_io_deq_bits_param;
	assign auto_in_d_bits_size = bundleIn_0_d_sink_io_deq_bits_size;
	assign auto_in_d_bits_source = bundleIn_0_d_sink_io_deq_bits_source;
	assign auto_in_d_bits_sink = bundleIn_0_d_sink_io_deq_bits_sink;
	assign auto_in_d_bits_denied = bundleIn_0_d_sink_io_deq_bits_denied;
	assign auto_in_d_bits_data = bundleIn_0_d_sink_io_deq_bits_data;
	assign auto_in_d_bits_corrupt = bundleIn_0_d_sink_io_deq_bits_corrupt;
	assign auto_out_a_mem_0_opcode = bundleOut_0_a_source_io_async_mem_0_opcode;
	assign auto_out_a_mem_0_address = bundleOut_0_a_source_io_async_mem_0_address;
	assign auto_out_a_mem_0_data = bundleOut_0_a_source_io_async_mem_0_data;
	assign auto_out_a_widx = bundleOut_0_a_source_io_async_widx;
	assign auto_out_a_safe_widx_valid = bundleOut_0_a_source_io_async_safe_widx_valid;
	assign auto_out_a_safe_source_reset_n = bundleOut_0_a_source_io_async_safe_source_reset_n;
	assign auto_out_d_ridx = bundleIn_0_d_sink_io_async_ridx;
	assign auto_out_d_safe_ridx_valid = bundleIn_0_d_sink_io_async_safe_ridx_valid;
	assign auto_out_d_safe_sink_reset_n = bundleIn_0_d_sink_io_async_safe_sink_reset_n;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = bundleOut_0_a_source_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = bundleIn_0_d_sink_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = bundleIn_0_d_sink_io_deq_bits_opcode;
	assign monitor_io_in_d_bits_param = bundleIn_0_d_sink_io_deq_bits_param;
	assign monitor_io_in_d_bits_size = bundleIn_0_d_sink_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = bundleIn_0_d_sink_io_deq_bits_source;
	assign monitor_io_in_d_bits_sink = bundleIn_0_d_sink_io_deq_bits_sink;
	assign monitor_io_in_d_bits_denied = bundleIn_0_d_sink_io_deq_bits_denied;
	assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_sink_io_deq_bits_corrupt;
	assign bundleOut_0_a_source_clock = clock;
	assign bundleOut_0_a_source_reset = reset;
	assign bundleOut_0_a_source_io_enq_valid = auto_in_a_valid;
	assign bundleOut_0_a_source_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign bundleOut_0_a_source_io_enq_bits_address = auto_in_a_bits_address;
	assign bundleOut_0_a_source_io_enq_bits_data = auto_in_a_bits_data;
	assign bundleOut_0_a_source_io_async_ridx = auto_out_a_ridx;
	assign bundleOut_0_a_source_io_async_safe_ridx_valid = auto_out_a_safe_ridx_valid;
	assign bundleOut_0_a_source_io_async_safe_sink_reset_n = auto_out_a_safe_sink_reset_n;
	assign bundleIn_0_d_sink_clock = clock;
	assign bundleIn_0_d_sink_reset = reset;
	assign bundleIn_0_d_sink_io_deq_ready = auto_in_d_ready;
	assign bundleIn_0_d_sink_io_async_mem_0_opcode = auto_out_d_mem_0_opcode;
	assign bundleIn_0_d_sink_io_async_mem_0_size = auto_out_d_mem_0_size;
	assign bundleIn_0_d_sink_io_async_mem_0_source = auto_out_d_mem_0_source;
	assign bundleIn_0_d_sink_io_async_mem_0_data = auto_out_d_mem_0_data;
	assign bundleIn_0_d_sink_io_async_widx = auto_out_d_widx;
	assign bundleIn_0_d_sink_io_async_safe_widx_valid = auto_out_d_safe_widx_valid;
	assign bundleIn_0_d_sink_io_async_safe_source_reset_n = auto_out_d_safe_source_reset_n;
endmodule
module AsyncQueueSource_1 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_resumereq,
	io_enq_bits_ackhavereset,
	io_enq_bits_hrmask_0,
	io_async_mem_0_resumereq,
	io_async_mem_0_ackhavereset,
	io_async_mem_0_hrmask_0,
	io_async_ridx,
	io_async_widx,
	io_async_safe_ridx_valid,
	io_async_safe_widx_valid,
	io_async_safe_source_reset_n,
	io_async_safe_sink_reset_n
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input io_enq_bits_resumereq;
	input io_enq_bits_ackhavereset;
	input io_enq_bits_hrmask_0;
	output wire io_async_mem_0_resumereq;
	output wire io_async_mem_0_ackhavereset;
	output wire io_async_mem_0_hrmask_0;
	input io_async_ridx;
	output wire io_async_widx;
	input io_async_safe_ridx_valid;
	output wire io_async_safe_widx_valid;
	output wire io_async_safe_source_reset_n;
	input io_async_safe_sink_reset_n;
	wire ridx_ridx_gray_clock;
	wire ridx_ridx_gray_reset;
	wire ridx_ridx_gray_io_d;
	wire ridx_ridx_gray_io_q;
	wire source_valid_0_io_in;
	wire source_valid_0_io_out;
	wire source_valid_0_clock;
	wire source_valid_0_reset;
	wire source_valid_1_io_in;
	wire source_valid_1_io_out;
	wire source_valid_1_clock;
	wire source_valid_1_reset;
	wire sink_extend_io_in;
	wire sink_extend_io_out;
	wire sink_extend_clock;
	wire sink_extend_reset;
	wire sink_valid_io_in;
	wire sink_valid_io_out;
	wire sink_valid_clock;
	wire sink_valid_reset;
	reg mem_0_resumereq;
	reg mem_0_ackhavereset;
	reg mem_0_hrmask_0;
	wire _widx_T_1 = io_enq_ready & io_enq_valid;
	wire sink_ready = sink_valid_io_out;
	wire _widx_T_2 = ~sink_ready;
	reg widx_widx_bin;
	wire widx_incremented = (_widx_T_2 ? 1'h0 : widx_widx_bin + _widx_T_1);
	wire ridx = ridx_ridx_gray_io_q;
	reg ready_reg;
	reg widx_gray;
	AsyncResetSynchronizerShiftReg_w1_d3_i0 ridx_ridx_gray(
		.clock(ridx_ridx_gray_clock),
		.reset(ridx_ridx_gray_reset),
		.io_d(ridx_ridx_gray_io_d),
		.io_q(ridx_ridx_gray_io_q)
	);
	AsyncValidSync source_valid_0(
		.io_in(source_valid_0_io_in),
		.io_out(source_valid_0_io_out),
		.clock(source_valid_0_clock),
		.reset(source_valid_0_reset)
	);
	AsyncValidSync source_valid_1(
		.io_in(source_valid_1_io_in),
		.io_out(source_valid_1_io_out),
		.clock(source_valid_1_clock),
		.reset(source_valid_1_reset)
	);
	AsyncValidSync sink_extend(
		.io_in(sink_extend_io_in),
		.io_out(sink_extend_io_out),
		.clock(sink_extend_clock),
		.reset(sink_extend_reset)
	);
	AsyncValidSync sink_valid(
		.io_in(sink_valid_io_in),
		.io_out(sink_valid_io_out),
		.clock(sink_valid_clock),
		.reset(sink_valid_reset)
	);
	assign io_enq_ready = ready_reg & sink_ready;
	assign io_async_mem_0_resumereq = mem_0_resumereq;
	assign io_async_mem_0_ackhavereset = mem_0_ackhavereset;
	assign io_async_mem_0_hrmask_0 = mem_0_hrmask_0;
	assign io_async_widx = widx_gray;
	assign io_async_safe_widx_valid = source_valid_1_io_out;
	assign io_async_safe_source_reset_n = ~reset;
	assign ridx_ridx_gray_clock = clock;
	assign ridx_ridx_gray_reset = reset;
	assign ridx_ridx_gray_io_d = io_async_ridx;
	assign source_valid_0_io_in = 1'h1;
	assign source_valid_0_clock = clock;
	assign source_valid_0_reset = reset | ~io_async_safe_sink_reset_n;
	assign source_valid_1_io_in = source_valid_0_io_out;
	assign source_valid_1_clock = clock;
	assign source_valid_1_reset = reset | ~io_async_safe_sink_reset_n;
	assign sink_extend_io_in = io_async_safe_ridx_valid;
	assign sink_extend_clock = clock;
	assign sink_extend_reset = reset | ~io_async_safe_sink_reset_n;
	assign sink_valid_io_in = sink_extend_io_out;
	assign sink_valid_clock = clock;
	assign sink_valid_reset = reset;
	always @(posedge clock) begin
		if (_widx_T_1)
			mem_0_resumereq <= io_enq_bits_resumereq;
		if (_widx_T_1)
			mem_0_ackhavereset <= io_enq_bits_ackhavereset;
		if (_widx_T_1)
			mem_0_hrmask_0 <= io_enq_bits_hrmask_0;
	end
	always @(posedge clock or posedge reset)
		if (reset)
			widx_widx_bin <= 1'h0;
		else if (_widx_T_2)
			widx_widx_bin <= 1'h0;
		else
			widx_widx_bin <= widx_widx_bin + _widx_T_1;
	always @(posedge clock or posedge reset)
		if (reset)
			ready_reg <= 1'h0;
		else
			ready_reg <= sink_ready & (widx_incremented != (ridx ^ 1'h1));
	always @(posedge clock or posedge reset)
		if (reset)
			widx_gray <= 1'h0;
		else if (_widx_T_2)
			widx_gray <= 1'h0;
		else
			widx_gray <= widx_widx_bin + _widx_T_1;
endmodule
module TLDebugModuleOuterAsync (
	auto_asource_out_a_mem_0_opcode,
	auto_asource_out_a_mem_0_address,
	auto_asource_out_a_mem_0_data,
	auto_asource_out_a_ridx,
	auto_asource_out_a_widx,
	auto_asource_out_a_safe_ridx_valid,
	auto_asource_out_a_safe_widx_valid,
	auto_asource_out_a_safe_source_reset_n,
	auto_asource_out_a_safe_sink_reset_n,
	auto_asource_out_d_mem_0_opcode,
	auto_asource_out_d_mem_0_size,
	auto_asource_out_d_mem_0_source,
	auto_asource_out_d_mem_0_data,
	auto_asource_out_d_ridx,
	auto_asource_out_d_widx,
	auto_asource_out_d_safe_ridx_valid,
	auto_asource_out_d_safe_widx_valid,
	auto_asource_out_d_safe_source_reset_n,
	auto_asource_out_d_safe_sink_reset_n,
	auto_intsource_out_sync_0,
	io_dmi_clock,
	io_dmi_reset,
	io_dmi_req_ready,
	io_dmi_req_valid,
	io_dmi_req_bits_addr,
	io_dmi_req_bits_data,
	io_dmi_req_bits_op,
	io_dmi_resp_ready,
	io_dmi_resp_valid,
	io_dmi_resp_bits_data,
	io_dmi_resp_bits_resp,
	io_ctrl_dmactive,
	io_ctrl_dmactiveAck,
	io_innerCtrl_mem_0_resumereq,
	io_innerCtrl_mem_0_ackhavereset,
	io_innerCtrl_mem_0_hrmask_0,
	io_innerCtrl_ridx,
	io_innerCtrl_widx,
	io_innerCtrl_safe_ridx_valid,
	io_innerCtrl_safe_widx_valid,
	io_innerCtrl_safe_source_reset_n,
	io_innerCtrl_safe_sink_reset_n,
	io_hgDebugInt_0
);
	output wire [2:0] auto_asource_out_a_mem_0_opcode;
	output wire [8:0] auto_asource_out_a_mem_0_address;
	output wire [31:0] auto_asource_out_a_mem_0_data;
	input auto_asource_out_a_ridx;
	output wire auto_asource_out_a_widx;
	input auto_asource_out_a_safe_ridx_valid;
	output wire auto_asource_out_a_safe_widx_valid;
	output wire auto_asource_out_a_safe_source_reset_n;
	input auto_asource_out_a_safe_sink_reset_n;
	input [2:0] auto_asource_out_d_mem_0_opcode;
	input [1:0] auto_asource_out_d_mem_0_size;
	input auto_asource_out_d_mem_0_source;
	input [31:0] auto_asource_out_d_mem_0_data;
	output wire auto_asource_out_d_ridx;
	input auto_asource_out_d_widx;
	output wire auto_asource_out_d_safe_ridx_valid;
	input auto_asource_out_d_safe_widx_valid;
	input auto_asource_out_d_safe_source_reset_n;
	output wire auto_asource_out_d_safe_sink_reset_n;
	output wire auto_intsource_out_sync_0;
	input io_dmi_clock;
	input io_dmi_reset;
	output wire io_dmi_req_ready;
	input io_dmi_req_valid;
	input [6:0] io_dmi_req_bits_addr;
	input [31:0] io_dmi_req_bits_data;
	input [1:0] io_dmi_req_bits_op;
	input io_dmi_resp_ready;
	output wire io_dmi_resp_valid;
	output wire [31:0] io_dmi_resp_bits_data;
	output wire [1:0] io_dmi_resp_bits_resp;
	output wire io_ctrl_dmactive;
	input io_ctrl_dmactiveAck;
	output wire io_innerCtrl_mem_0_resumereq;
	output wire io_innerCtrl_mem_0_ackhavereset;
	output wire io_innerCtrl_mem_0_hrmask_0;
	input io_innerCtrl_ridx;
	output wire io_innerCtrl_widx;
	input io_innerCtrl_safe_ridx_valid;
	output wire io_innerCtrl_safe_widx_valid;
	output wire io_innerCtrl_safe_source_reset_n;
	input io_innerCtrl_safe_sink_reset_n;
	input io_hgDebugInt_0;
	wire dmiXbar_clock;
	wire dmiXbar_reset;
	wire dmiXbar_auto_in_a_ready;
	wire dmiXbar_auto_in_a_valid;
	wire [2:0] dmiXbar_auto_in_a_bits_opcode;
	wire [8:0] dmiXbar_auto_in_a_bits_address;
	wire [31:0] dmiXbar_auto_in_a_bits_data;
	wire dmiXbar_auto_in_d_ready;
	wire dmiXbar_auto_in_d_valid;
	wire dmiXbar_auto_in_d_bits_denied;
	wire [31:0] dmiXbar_auto_in_d_bits_data;
	wire dmiXbar_auto_in_d_bits_corrupt;
	wire dmiXbar_auto_out_1_a_ready;
	wire dmiXbar_auto_out_1_a_valid;
	wire [2:0] dmiXbar_auto_out_1_a_bits_opcode;
	wire [6:0] dmiXbar_auto_out_1_a_bits_address;
	wire [31:0] dmiXbar_auto_out_1_a_bits_data;
	wire dmiXbar_auto_out_1_d_ready;
	wire dmiXbar_auto_out_1_d_valid;
	wire [2:0] dmiXbar_auto_out_1_d_bits_opcode;
	wire [31:0] dmiXbar_auto_out_1_d_bits_data;
	wire dmiXbar_auto_out_0_a_ready;
	wire dmiXbar_auto_out_0_a_valid;
	wire [2:0] dmiXbar_auto_out_0_a_bits_opcode;
	wire [8:0] dmiXbar_auto_out_0_a_bits_address;
	wire [31:0] dmiXbar_auto_out_0_a_bits_data;
	wire dmiXbar_auto_out_0_d_ready;
	wire dmiXbar_auto_out_0_d_valid;
	wire [2:0] dmiXbar_auto_out_0_d_bits_opcode;
	wire [1:0] dmiXbar_auto_out_0_d_bits_param;
	wire [1:0] dmiXbar_auto_out_0_d_bits_size;
	wire dmiXbar_auto_out_0_d_bits_sink;
	wire dmiXbar_auto_out_0_d_bits_denied;
	wire [31:0] dmiXbar_auto_out_0_d_bits_data;
	wire dmiXbar_auto_out_0_d_bits_corrupt;
	wire dmi2tl_auto_out_a_ready;
	wire dmi2tl_auto_out_a_valid;
	wire [2:0] dmi2tl_auto_out_a_bits_opcode;
	wire [8:0] dmi2tl_auto_out_a_bits_address;
	wire [31:0] dmi2tl_auto_out_a_bits_data;
	wire dmi2tl_auto_out_d_ready;
	wire dmi2tl_auto_out_d_valid;
	wire dmi2tl_auto_out_d_bits_denied;
	wire [31:0] dmi2tl_auto_out_d_bits_data;
	wire dmi2tl_auto_out_d_bits_corrupt;
	wire dmi2tl_io_dmi_req_ready;
	wire dmi2tl_io_dmi_req_valid;
	wire [6:0] dmi2tl_io_dmi_req_bits_addr;
	wire [31:0] dmi2tl_io_dmi_req_bits_data;
	wire [1:0] dmi2tl_io_dmi_req_bits_op;
	wire dmi2tl_io_dmi_resp_ready;
	wire dmi2tl_io_dmi_resp_valid;
	wire [31:0] dmi2tl_io_dmi_resp_bits_data;
	wire [1:0] dmi2tl_io_dmi_resp_bits_resp;
	wire dmOuter_clock;
	wire dmOuter_reset;
	wire dmOuter_auto_dmi_in_a_ready;
	wire dmOuter_auto_dmi_in_a_valid;
	wire [2:0] dmOuter_auto_dmi_in_a_bits_opcode;
	wire [6:0] dmOuter_auto_dmi_in_a_bits_address;
	wire [31:0] dmOuter_auto_dmi_in_a_bits_data;
	wire dmOuter_auto_dmi_in_d_ready;
	wire dmOuter_auto_dmi_in_d_valid;
	wire [2:0] dmOuter_auto_dmi_in_d_bits_opcode;
	wire [31:0] dmOuter_auto_dmi_in_d_bits_data;
	wire dmOuter_auto_int_out_0;
	wire dmOuter_io_ctrl_dmactive;
	wire dmOuter_io_ctrl_dmactiveAck;
	wire dmOuter_io_innerCtrl_ready;
	wire dmOuter_io_innerCtrl_valid;
	wire dmOuter_io_innerCtrl_bits_resumereq;
	wire [9:0] dmOuter_io_innerCtrl_bits_hartsel;
	wire dmOuter_io_innerCtrl_bits_ackhavereset;
	wire dmOuter_io_innerCtrl_bits_hrmask_0;
	wire dmOuter_io_hgDebugInt_0;
	wire intsource_auto_in_0;
	wire intsource_auto_out_sync_0;
	wire dmiBypass_clock;
	wire dmiBypass_reset;
	wire dmiBypass_auto_node_out_out_a_ready;
	wire dmiBypass_auto_node_out_out_a_valid;
	wire [2:0] dmiBypass_auto_node_out_out_a_bits_opcode;
	wire [8:0] dmiBypass_auto_node_out_out_a_bits_address;
	wire [31:0] dmiBypass_auto_node_out_out_a_bits_data;
	wire dmiBypass_auto_node_out_out_d_ready;
	wire dmiBypass_auto_node_out_out_d_valid;
	wire [2:0] dmiBypass_auto_node_out_out_d_bits_opcode;
	wire [1:0] dmiBypass_auto_node_out_out_d_bits_param;
	wire [1:0] dmiBypass_auto_node_out_out_d_bits_size;
	wire dmiBypass_auto_node_out_out_d_bits_source;
	wire dmiBypass_auto_node_out_out_d_bits_sink;
	wire dmiBypass_auto_node_out_out_d_bits_denied;
	wire [31:0] dmiBypass_auto_node_out_out_d_bits_data;
	wire dmiBypass_auto_node_out_out_d_bits_corrupt;
	wire dmiBypass_auto_node_in_in_a_ready;
	wire dmiBypass_auto_node_in_in_a_valid;
	wire [2:0] dmiBypass_auto_node_in_in_a_bits_opcode;
	wire [8:0] dmiBypass_auto_node_in_in_a_bits_address;
	wire [31:0] dmiBypass_auto_node_in_in_a_bits_data;
	wire dmiBypass_auto_node_in_in_d_ready;
	wire dmiBypass_auto_node_in_in_d_valid;
	wire [2:0] dmiBypass_auto_node_in_in_d_bits_opcode;
	wire [1:0] dmiBypass_auto_node_in_in_d_bits_param;
	wire [1:0] dmiBypass_auto_node_in_in_d_bits_size;
	wire dmiBypass_auto_node_in_in_d_bits_sink;
	wire dmiBypass_auto_node_in_in_d_bits_denied;
	wire [31:0] dmiBypass_auto_node_in_in_d_bits_data;
	wire dmiBypass_auto_node_in_in_d_bits_corrupt;
	wire dmiBypass_io_bypass;
	wire asource_clock;
	wire asource_reset;
	wire asource_auto_in_a_ready;
	wire asource_auto_in_a_valid;
	wire [2:0] asource_auto_in_a_bits_opcode;
	wire [8:0] asource_auto_in_a_bits_address;
	wire [31:0] asource_auto_in_a_bits_data;
	wire asource_auto_in_d_ready;
	wire asource_auto_in_d_valid;
	wire [2:0] asource_auto_in_d_bits_opcode;
	wire [1:0] asource_auto_in_d_bits_param;
	wire [1:0] asource_auto_in_d_bits_size;
	wire asource_auto_in_d_bits_source;
	wire asource_auto_in_d_bits_sink;
	wire asource_auto_in_d_bits_denied;
	wire [31:0] asource_auto_in_d_bits_data;
	wire asource_auto_in_d_bits_corrupt;
	wire [2:0] asource_auto_out_a_mem_0_opcode;
	wire [8:0] asource_auto_out_a_mem_0_address;
	wire [31:0] asource_auto_out_a_mem_0_data;
	wire asource_auto_out_a_ridx;
	wire asource_auto_out_a_widx;
	wire asource_auto_out_a_safe_ridx_valid;
	wire asource_auto_out_a_safe_widx_valid;
	wire asource_auto_out_a_safe_source_reset_n;
	wire asource_auto_out_a_safe_sink_reset_n;
	wire [2:0] asource_auto_out_d_mem_0_opcode;
	wire [1:0] asource_auto_out_d_mem_0_size;
	wire asource_auto_out_d_mem_0_source;
	wire [31:0] asource_auto_out_d_mem_0_data;
	wire asource_auto_out_d_ridx;
	wire asource_auto_out_d_widx;
	wire asource_auto_out_d_safe_ridx_valid;
	wire asource_auto_out_d_safe_widx_valid;
	wire asource_auto_out_d_safe_source_reset_n;
	wire asource_auto_out_d_safe_sink_reset_n;
	wire dmactiveAck_dmactiveAckSync_clock;
	wire dmactiveAck_dmactiveAckSync_reset;
	wire dmactiveAck_dmactiveAckSync_io_d;
	wire dmactiveAck_dmactiveAckSync_io_q;
	wire io_innerCtrl_source_clock;
	wire io_innerCtrl_source_reset;
	wire io_innerCtrl_source_io_enq_ready;
	wire io_innerCtrl_source_io_enq_valid;
	wire io_innerCtrl_source_io_enq_bits_resumereq;
	wire io_innerCtrl_source_io_enq_bits_ackhavereset;
	wire io_innerCtrl_source_io_enq_bits_hrmask_0;
	wire io_innerCtrl_source_io_async_mem_0_resumereq;
	wire io_innerCtrl_source_io_async_mem_0_ackhavereset;
	wire io_innerCtrl_source_io_async_mem_0_hrmask_0;
	wire io_innerCtrl_source_io_async_ridx;
	wire io_innerCtrl_source_io_async_widx;
	wire io_innerCtrl_source_io_async_safe_ridx_valid;
	wire io_innerCtrl_source_io_async_safe_widx_valid;
	wire io_innerCtrl_source_io_async_safe_source_reset_n;
	wire io_innerCtrl_source_io_async_safe_sink_reset_n;
	wire dmactiveAck = dmactiveAck_dmactiveAckSync_io_q;
	TLXbar_8 dmiXbar(
		.clock(dmiXbar_clock),
		.reset(dmiXbar_reset),
		.auto_in_a_ready(dmiXbar_auto_in_a_ready),
		.auto_in_a_valid(dmiXbar_auto_in_a_valid),
		.auto_in_a_bits_opcode(dmiXbar_auto_in_a_bits_opcode),
		.auto_in_a_bits_address(dmiXbar_auto_in_a_bits_address),
		.auto_in_a_bits_data(dmiXbar_auto_in_a_bits_data),
		.auto_in_d_ready(dmiXbar_auto_in_d_ready),
		.auto_in_d_valid(dmiXbar_auto_in_d_valid),
		.auto_in_d_bits_denied(dmiXbar_auto_in_d_bits_denied),
		.auto_in_d_bits_data(dmiXbar_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(dmiXbar_auto_in_d_bits_corrupt),
		.auto_out_1_a_ready(dmiXbar_auto_out_1_a_ready),
		.auto_out_1_a_valid(dmiXbar_auto_out_1_a_valid),
		.auto_out_1_a_bits_opcode(dmiXbar_auto_out_1_a_bits_opcode),
		.auto_out_1_a_bits_address(dmiXbar_auto_out_1_a_bits_address),
		.auto_out_1_a_bits_data(dmiXbar_auto_out_1_a_bits_data),
		.auto_out_1_d_ready(dmiXbar_auto_out_1_d_ready),
		.auto_out_1_d_valid(dmiXbar_auto_out_1_d_valid),
		.auto_out_1_d_bits_opcode(dmiXbar_auto_out_1_d_bits_opcode),
		.auto_out_1_d_bits_data(dmiXbar_auto_out_1_d_bits_data),
		.auto_out_0_a_ready(dmiXbar_auto_out_0_a_ready),
		.auto_out_0_a_valid(dmiXbar_auto_out_0_a_valid),
		.auto_out_0_a_bits_opcode(dmiXbar_auto_out_0_a_bits_opcode),
		.auto_out_0_a_bits_address(dmiXbar_auto_out_0_a_bits_address),
		.auto_out_0_a_bits_data(dmiXbar_auto_out_0_a_bits_data),
		.auto_out_0_d_ready(dmiXbar_auto_out_0_d_ready),
		.auto_out_0_d_valid(dmiXbar_auto_out_0_d_valid),
		.auto_out_0_d_bits_opcode(dmiXbar_auto_out_0_d_bits_opcode),
		.auto_out_0_d_bits_param(dmiXbar_auto_out_0_d_bits_param),
		.auto_out_0_d_bits_size(dmiXbar_auto_out_0_d_bits_size),
		.auto_out_0_d_bits_sink(dmiXbar_auto_out_0_d_bits_sink),
		.auto_out_0_d_bits_denied(dmiXbar_auto_out_0_d_bits_denied),
		.auto_out_0_d_bits_data(dmiXbar_auto_out_0_d_bits_data),
		.auto_out_0_d_bits_corrupt(dmiXbar_auto_out_0_d_bits_corrupt)
	);
	DMIToTL dmi2tl(
		.auto_out_a_ready(dmi2tl_auto_out_a_ready),
		.auto_out_a_valid(dmi2tl_auto_out_a_valid),
		.auto_out_a_bits_opcode(dmi2tl_auto_out_a_bits_opcode),
		.auto_out_a_bits_address(dmi2tl_auto_out_a_bits_address),
		.auto_out_a_bits_data(dmi2tl_auto_out_a_bits_data),
		.auto_out_d_ready(dmi2tl_auto_out_d_ready),
		.auto_out_d_valid(dmi2tl_auto_out_d_valid),
		.auto_out_d_bits_denied(dmi2tl_auto_out_d_bits_denied),
		.auto_out_d_bits_data(dmi2tl_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(dmi2tl_auto_out_d_bits_corrupt),
		.io_dmi_req_ready(dmi2tl_io_dmi_req_ready),
		.io_dmi_req_valid(dmi2tl_io_dmi_req_valid),
		.io_dmi_req_bits_addr(dmi2tl_io_dmi_req_bits_addr),
		.io_dmi_req_bits_data(dmi2tl_io_dmi_req_bits_data),
		.io_dmi_req_bits_op(dmi2tl_io_dmi_req_bits_op),
		.io_dmi_resp_ready(dmi2tl_io_dmi_resp_ready),
		.io_dmi_resp_valid(dmi2tl_io_dmi_resp_valid),
		.io_dmi_resp_bits_data(dmi2tl_io_dmi_resp_bits_data),
		.io_dmi_resp_bits_resp(dmi2tl_io_dmi_resp_bits_resp)
	);
	TLDebugModuleOuter dmOuter(
		.clock(dmOuter_clock),
		.reset(dmOuter_reset),
		.auto_dmi_in_a_ready(dmOuter_auto_dmi_in_a_ready),
		.auto_dmi_in_a_valid(dmOuter_auto_dmi_in_a_valid),
		.auto_dmi_in_a_bits_opcode(dmOuter_auto_dmi_in_a_bits_opcode),
		.auto_dmi_in_a_bits_address(dmOuter_auto_dmi_in_a_bits_address),
		.auto_dmi_in_a_bits_data(dmOuter_auto_dmi_in_a_bits_data),
		.auto_dmi_in_d_ready(dmOuter_auto_dmi_in_d_ready),
		.auto_dmi_in_d_valid(dmOuter_auto_dmi_in_d_valid),
		.auto_dmi_in_d_bits_opcode(dmOuter_auto_dmi_in_d_bits_opcode),
		.auto_dmi_in_d_bits_data(dmOuter_auto_dmi_in_d_bits_data),
		.auto_int_out_0(dmOuter_auto_int_out_0),
		.io_ctrl_dmactive(dmOuter_io_ctrl_dmactive),
		.io_ctrl_dmactiveAck(dmOuter_io_ctrl_dmactiveAck),
		.io_innerCtrl_ready(dmOuter_io_innerCtrl_ready),
		.io_innerCtrl_valid(dmOuter_io_innerCtrl_valid),
		.io_innerCtrl_bits_resumereq(dmOuter_io_innerCtrl_bits_resumereq),
		.io_innerCtrl_bits_hartsel(dmOuter_io_innerCtrl_bits_hartsel),
		.io_innerCtrl_bits_ackhavereset(dmOuter_io_innerCtrl_bits_ackhavereset),
		.io_innerCtrl_bits_hrmask_0(dmOuter_io_innerCtrl_bits_hrmask_0),
		.io_hgDebugInt_0(dmOuter_io_hgDebugInt_0)
	);
	IntSyncCrossingSource_4 intsource(
		.auto_in_0(intsource_auto_in_0),
		.auto_out_sync_0(intsource_auto_out_sync_0)
	);
	TLBusBypass dmiBypass(
		.clock(dmiBypass_clock),
		.reset(dmiBypass_reset),
		.auto_node_out_out_a_ready(dmiBypass_auto_node_out_out_a_ready),
		.auto_node_out_out_a_valid(dmiBypass_auto_node_out_out_a_valid),
		.auto_node_out_out_a_bits_opcode(dmiBypass_auto_node_out_out_a_bits_opcode),
		.auto_node_out_out_a_bits_address(dmiBypass_auto_node_out_out_a_bits_address),
		.auto_node_out_out_a_bits_data(dmiBypass_auto_node_out_out_a_bits_data),
		.auto_node_out_out_d_ready(dmiBypass_auto_node_out_out_d_ready),
		.auto_node_out_out_d_valid(dmiBypass_auto_node_out_out_d_valid),
		.auto_node_out_out_d_bits_opcode(dmiBypass_auto_node_out_out_d_bits_opcode),
		.auto_node_out_out_d_bits_param(dmiBypass_auto_node_out_out_d_bits_param),
		.auto_node_out_out_d_bits_size(dmiBypass_auto_node_out_out_d_bits_size),
		.auto_node_out_out_d_bits_source(dmiBypass_auto_node_out_out_d_bits_source),
		.auto_node_out_out_d_bits_sink(dmiBypass_auto_node_out_out_d_bits_sink),
		.auto_node_out_out_d_bits_denied(dmiBypass_auto_node_out_out_d_bits_denied),
		.auto_node_out_out_d_bits_data(dmiBypass_auto_node_out_out_d_bits_data),
		.auto_node_out_out_d_bits_corrupt(dmiBypass_auto_node_out_out_d_bits_corrupt),
		.auto_node_in_in_a_ready(dmiBypass_auto_node_in_in_a_ready),
		.auto_node_in_in_a_valid(dmiBypass_auto_node_in_in_a_valid),
		.auto_node_in_in_a_bits_opcode(dmiBypass_auto_node_in_in_a_bits_opcode),
		.auto_node_in_in_a_bits_address(dmiBypass_auto_node_in_in_a_bits_address),
		.auto_node_in_in_a_bits_data(dmiBypass_auto_node_in_in_a_bits_data),
		.auto_node_in_in_d_ready(dmiBypass_auto_node_in_in_d_ready),
		.auto_node_in_in_d_valid(dmiBypass_auto_node_in_in_d_valid),
		.auto_node_in_in_d_bits_opcode(dmiBypass_auto_node_in_in_d_bits_opcode),
		.auto_node_in_in_d_bits_param(dmiBypass_auto_node_in_in_d_bits_param),
		.auto_node_in_in_d_bits_size(dmiBypass_auto_node_in_in_d_bits_size),
		.auto_node_in_in_d_bits_sink(dmiBypass_auto_node_in_in_d_bits_sink),
		.auto_node_in_in_d_bits_denied(dmiBypass_auto_node_in_in_d_bits_denied),
		.auto_node_in_in_d_bits_data(dmiBypass_auto_node_in_in_d_bits_data),
		.auto_node_in_in_d_bits_corrupt(dmiBypass_auto_node_in_in_d_bits_corrupt),
		.io_bypass(dmiBypass_io_bypass)
	);
	TLAsyncCrossingSource asource(
		.clock(asource_clock),
		.reset(asource_reset),
		.auto_in_a_ready(asource_auto_in_a_ready),
		.auto_in_a_valid(asource_auto_in_a_valid),
		.auto_in_a_bits_opcode(asource_auto_in_a_bits_opcode),
		.auto_in_a_bits_address(asource_auto_in_a_bits_address),
		.auto_in_a_bits_data(asource_auto_in_a_bits_data),
		.auto_in_d_ready(asource_auto_in_d_ready),
		.auto_in_d_valid(asource_auto_in_d_valid),
		.auto_in_d_bits_opcode(asource_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(asource_auto_in_d_bits_param),
		.auto_in_d_bits_size(asource_auto_in_d_bits_size),
		.auto_in_d_bits_source(asource_auto_in_d_bits_source),
		.auto_in_d_bits_sink(asource_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(asource_auto_in_d_bits_denied),
		.auto_in_d_bits_data(asource_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(asource_auto_in_d_bits_corrupt),
		.auto_out_a_mem_0_opcode(asource_auto_out_a_mem_0_opcode),
		.auto_out_a_mem_0_address(asource_auto_out_a_mem_0_address),
		.auto_out_a_mem_0_data(asource_auto_out_a_mem_0_data),
		.auto_out_a_ridx(asource_auto_out_a_ridx),
		.auto_out_a_widx(asource_auto_out_a_widx),
		.auto_out_a_safe_ridx_valid(asource_auto_out_a_safe_ridx_valid),
		.auto_out_a_safe_widx_valid(asource_auto_out_a_safe_widx_valid),
		.auto_out_a_safe_source_reset_n(asource_auto_out_a_safe_source_reset_n),
		.auto_out_a_safe_sink_reset_n(asource_auto_out_a_safe_sink_reset_n),
		.auto_out_d_mem_0_opcode(asource_auto_out_d_mem_0_opcode),
		.auto_out_d_mem_0_size(asource_auto_out_d_mem_0_size),
		.auto_out_d_mem_0_source(asource_auto_out_d_mem_0_source),
		.auto_out_d_mem_0_data(asource_auto_out_d_mem_0_data),
		.auto_out_d_ridx(asource_auto_out_d_ridx),
		.auto_out_d_widx(asource_auto_out_d_widx),
		.auto_out_d_safe_ridx_valid(asource_auto_out_d_safe_ridx_valid),
		.auto_out_d_safe_widx_valid(asource_auto_out_d_safe_widx_valid),
		.auto_out_d_safe_source_reset_n(asource_auto_out_d_safe_source_reset_n),
		.auto_out_d_safe_sink_reset_n(asource_auto_out_d_safe_sink_reset_n)
	);
	AsyncResetSynchronizerShiftReg_w1_d3_i0 dmactiveAck_dmactiveAckSync(
		.clock(dmactiveAck_dmactiveAckSync_clock),
		.reset(dmactiveAck_dmactiveAckSync_reset),
		.io_d(dmactiveAck_dmactiveAckSync_io_d),
		.io_q(dmactiveAck_dmactiveAckSync_io_q)
	);
	AsyncQueueSource_1 io_innerCtrl_source(
		.clock(io_innerCtrl_source_clock),
		.reset(io_innerCtrl_source_reset),
		.io_enq_ready(io_innerCtrl_source_io_enq_ready),
		.io_enq_valid(io_innerCtrl_source_io_enq_valid),
		.io_enq_bits_resumereq(io_innerCtrl_source_io_enq_bits_resumereq),
		.io_enq_bits_ackhavereset(io_innerCtrl_source_io_enq_bits_ackhavereset),
		.io_enq_bits_hrmask_0(io_innerCtrl_source_io_enq_bits_hrmask_0),
		.io_async_mem_0_resumereq(io_innerCtrl_source_io_async_mem_0_resumereq),
		.io_async_mem_0_ackhavereset(io_innerCtrl_source_io_async_mem_0_ackhavereset),
		.io_async_mem_0_hrmask_0(io_innerCtrl_source_io_async_mem_0_hrmask_0),
		.io_async_ridx(io_innerCtrl_source_io_async_ridx),
		.io_async_widx(io_innerCtrl_source_io_async_widx),
		.io_async_safe_ridx_valid(io_innerCtrl_source_io_async_safe_ridx_valid),
		.io_async_safe_widx_valid(io_innerCtrl_source_io_async_safe_widx_valid),
		.io_async_safe_source_reset_n(io_innerCtrl_source_io_async_safe_source_reset_n),
		.io_async_safe_sink_reset_n(io_innerCtrl_source_io_async_safe_sink_reset_n)
	);
	assign auto_asource_out_a_mem_0_opcode = asource_auto_out_a_mem_0_opcode;
	assign auto_asource_out_a_mem_0_address = asource_auto_out_a_mem_0_address;
	assign auto_asource_out_a_mem_0_data = asource_auto_out_a_mem_0_data;
	assign auto_asource_out_a_widx = asource_auto_out_a_widx;
	assign auto_asource_out_a_safe_widx_valid = asource_auto_out_a_safe_widx_valid;
	assign auto_asource_out_a_safe_source_reset_n = asource_auto_out_a_safe_source_reset_n;
	assign auto_asource_out_d_ridx = asource_auto_out_d_ridx;
	assign auto_asource_out_d_safe_ridx_valid = asource_auto_out_d_safe_ridx_valid;
	assign auto_asource_out_d_safe_sink_reset_n = asource_auto_out_d_safe_sink_reset_n;
	assign auto_intsource_out_sync_0 = intsource_auto_out_sync_0;
	assign io_dmi_req_ready = dmi2tl_io_dmi_req_ready;
	assign io_dmi_resp_valid = dmi2tl_io_dmi_resp_valid;
	assign io_dmi_resp_bits_data = dmi2tl_io_dmi_resp_bits_data;
	assign io_dmi_resp_bits_resp = dmi2tl_io_dmi_resp_bits_resp;
	assign io_ctrl_dmactive = dmOuter_io_ctrl_dmactive;
	assign io_innerCtrl_mem_0_resumereq = io_innerCtrl_source_io_async_mem_0_resumereq;
	assign io_innerCtrl_mem_0_ackhavereset = io_innerCtrl_source_io_async_mem_0_ackhavereset;
	assign io_innerCtrl_mem_0_hrmask_0 = io_innerCtrl_source_io_async_mem_0_hrmask_0;
	assign io_innerCtrl_widx = io_innerCtrl_source_io_async_widx;
	assign io_innerCtrl_safe_widx_valid = io_innerCtrl_source_io_async_safe_widx_valid;
	assign io_innerCtrl_safe_source_reset_n = io_innerCtrl_source_io_async_safe_source_reset_n;
	assign dmiXbar_clock = io_dmi_clock;
	assign dmiXbar_reset = io_dmi_reset;
	assign dmiXbar_auto_in_a_valid = dmi2tl_auto_out_a_valid;
	assign dmiXbar_auto_in_a_bits_opcode = dmi2tl_auto_out_a_bits_opcode;
	assign dmiXbar_auto_in_a_bits_address = dmi2tl_auto_out_a_bits_address;
	assign dmiXbar_auto_in_a_bits_data = dmi2tl_auto_out_a_bits_data;
	assign dmiXbar_auto_in_d_ready = dmi2tl_auto_out_d_ready;
	assign dmiXbar_auto_out_1_a_ready = dmOuter_auto_dmi_in_a_ready;
	assign dmiXbar_auto_out_1_d_valid = dmOuter_auto_dmi_in_d_valid;
	assign dmiXbar_auto_out_1_d_bits_opcode = dmOuter_auto_dmi_in_d_bits_opcode;
	assign dmiXbar_auto_out_1_d_bits_data = dmOuter_auto_dmi_in_d_bits_data;
	assign dmiXbar_auto_out_0_a_ready = dmiBypass_auto_node_in_in_a_ready;
	assign dmiXbar_auto_out_0_d_valid = dmiBypass_auto_node_in_in_d_valid;
	assign dmiXbar_auto_out_0_d_bits_opcode = dmiBypass_auto_node_in_in_d_bits_opcode;
	assign dmiXbar_auto_out_0_d_bits_param = dmiBypass_auto_node_in_in_d_bits_param;
	assign dmiXbar_auto_out_0_d_bits_size = dmiBypass_auto_node_in_in_d_bits_size;
	assign dmiXbar_auto_out_0_d_bits_sink = dmiBypass_auto_node_in_in_d_bits_sink;
	assign dmiXbar_auto_out_0_d_bits_denied = dmiBypass_auto_node_in_in_d_bits_denied;
	assign dmiXbar_auto_out_0_d_bits_data = dmiBypass_auto_node_in_in_d_bits_data;
	assign dmiXbar_auto_out_0_d_bits_corrupt = dmiBypass_auto_node_in_in_d_bits_corrupt;
	assign dmi2tl_auto_out_a_ready = dmiXbar_auto_in_a_ready;
	assign dmi2tl_auto_out_d_valid = dmiXbar_auto_in_d_valid;
	assign dmi2tl_auto_out_d_bits_denied = dmiXbar_auto_in_d_bits_denied;
	assign dmi2tl_auto_out_d_bits_data = dmiXbar_auto_in_d_bits_data;
	assign dmi2tl_auto_out_d_bits_corrupt = dmiXbar_auto_in_d_bits_corrupt;
	assign dmi2tl_io_dmi_req_valid = io_dmi_req_valid;
	assign dmi2tl_io_dmi_req_bits_addr = io_dmi_req_bits_addr;
	assign dmi2tl_io_dmi_req_bits_data = io_dmi_req_bits_data;
	assign dmi2tl_io_dmi_req_bits_op = io_dmi_req_bits_op;
	assign dmi2tl_io_dmi_resp_ready = io_dmi_resp_ready;
	assign dmOuter_clock = io_dmi_clock;
	assign dmOuter_reset = io_dmi_reset;
	assign dmOuter_auto_dmi_in_a_valid = dmiXbar_auto_out_1_a_valid;
	assign dmOuter_auto_dmi_in_a_bits_opcode = dmiXbar_auto_out_1_a_bits_opcode;
	assign dmOuter_auto_dmi_in_a_bits_address = dmiXbar_auto_out_1_a_bits_address;
	assign dmOuter_auto_dmi_in_a_bits_data = dmiXbar_auto_out_1_a_bits_data;
	assign dmOuter_auto_dmi_in_d_ready = dmiXbar_auto_out_1_d_ready;
	assign dmOuter_io_ctrl_dmactiveAck = dmactiveAck_dmactiveAckSync_io_q;
	assign dmOuter_io_innerCtrl_ready = io_innerCtrl_source_io_enq_ready;
	assign dmOuter_io_hgDebugInt_0 = io_hgDebugInt_0;
	assign intsource_auto_in_0 = dmOuter_auto_int_out_0;
	assign dmiBypass_clock = io_dmi_clock;
	assign dmiBypass_reset = io_dmi_reset;
	assign dmiBypass_auto_node_out_out_a_ready = asource_auto_in_a_ready;
	assign dmiBypass_auto_node_out_out_d_valid = asource_auto_in_d_valid;
	assign dmiBypass_auto_node_out_out_d_bits_opcode = asource_auto_in_d_bits_opcode;
	assign dmiBypass_auto_node_out_out_d_bits_param = asource_auto_in_d_bits_param;
	assign dmiBypass_auto_node_out_out_d_bits_size = asource_auto_in_d_bits_size;
	assign dmiBypass_auto_node_out_out_d_bits_source = asource_auto_in_d_bits_source;
	assign dmiBypass_auto_node_out_out_d_bits_sink = asource_auto_in_d_bits_sink;
	assign dmiBypass_auto_node_out_out_d_bits_denied = asource_auto_in_d_bits_denied;
	assign dmiBypass_auto_node_out_out_d_bits_data = asource_auto_in_d_bits_data;
	assign dmiBypass_auto_node_out_out_d_bits_corrupt = asource_auto_in_d_bits_corrupt;
	assign dmiBypass_auto_node_in_in_a_valid = dmiXbar_auto_out_0_a_valid;
	assign dmiBypass_auto_node_in_in_a_bits_opcode = dmiXbar_auto_out_0_a_bits_opcode;
	assign dmiBypass_auto_node_in_in_a_bits_address = dmiXbar_auto_out_0_a_bits_address;
	assign dmiBypass_auto_node_in_in_a_bits_data = dmiXbar_auto_out_0_a_bits_data;
	assign dmiBypass_auto_node_in_in_d_ready = dmiXbar_auto_out_0_d_ready;
	assign dmiBypass_io_bypass = ~io_ctrl_dmactive | ~dmactiveAck;
	assign asource_clock = io_dmi_clock;
	assign asource_reset = io_dmi_reset;
	assign asource_auto_in_a_valid = dmiBypass_auto_node_out_out_a_valid;
	assign asource_auto_in_a_bits_opcode = dmiBypass_auto_node_out_out_a_bits_opcode;
	assign asource_auto_in_a_bits_address = dmiBypass_auto_node_out_out_a_bits_address;
	assign asource_auto_in_a_bits_data = dmiBypass_auto_node_out_out_a_bits_data;
	assign asource_auto_in_d_ready = dmiBypass_auto_node_out_out_d_ready;
	assign asource_auto_out_a_ridx = auto_asource_out_a_ridx;
	assign asource_auto_out_a_safe_ridx_valid = auto_asource_out_a_safe_ridx_valid;
	assign asource_auto_out_a_safe_sink_reset_n = auto_asource_out_a_safe_sink_reset_n;
	assign asource_auto_out_d_mem_0_opcode = auto_asource_out_d_mem_0_opcode;
	assign asource_auto_out_d_mem_0_size = auto_asource_out_d_mem_0_size;
	assign asource_auto_out_d_mem_0_source = auto_asource_out_d_mem_0_source;
	assign asource_auto_out_d_mem_0_data = auto_asource_out_d_mem_0_data;
	assign asource_auto_out_d_widx = auto_asource_out_d_widx;
	assign asource_auto_out_d_safe_widx_valid = auto_asource_out_d_safe_widx_valid;
	assign asource_auto_out_d_safe_source_reset_n = auto_asource_out_d_safe_source_reset_n;
	assign dmactiveAck_dmactiveAckSync_clock = io_dmi_clock;
	assign dmactiveAck_dmactiveAckSync_reset = io_dmi_reset;
	assign dmactiveAck_dmactiveAckSync_io_d = io_ctrl_dmactiveAck;
	assign io_innerCtrl_source_clock = io_dmi_clock;
	assign io_innerCtrl_source_reset = io_dmi_reset;
	assign io_innerCtrl_source_io_enq_valid = dmOuter_io_innerCtrl_valid;
	assign io_innerCtrl_source_io_enq_bits_resumereq = dmOuter_io_innerCtrl_bits_resumereq;
	assign io_innerCtrl_source_io_enq_bits_ackhavereset = dmOuter_io_innerCtrl_bits_ackhavereset;
	assign io_innerCtrl_source_io_enq_bits_hrmask_0 = dmOuter_io_innerCtrl_bits_hrmask_0;
	assign io_innerCtrl_source_io_async_ridx = io_innerCtrl_ridx;
	assign io_innerCtrl_source_io_async_safe_ridx_valid = io_innerCtrl_safe_ridx_valid;
	assign io_innerCtrl_source_io_async_safe_sink_reset_n = io_innerCtrl_safe_sink_reset_n;
endmodule
module TLMonitor_41 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [1:0] io_in_a_bits_size;
	input io_in_a_bits_source;
	input [8:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_size;
	input io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = ~io_in_a_bits_source;
	wire [4:0] _is_aligned_mask_T_1 = 5'h03 << io_in_a_bits_size;
	wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0];
	wire [8:0] _GEN_71 = {7'd0, is_aligned_mask};
	wire [8:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 9'h000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 2'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_5 = ~_source_ok_T;
	wire [9:0] _T_7 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_15 = io_in_a_bits_opcode == 3'h6;
	wire [9:0] _T_23 = $signed(_T_7) & -10'sh040;
	wire _T_24 = $signed(_T_23) == 10'sh000;
	wire [8:0] _T_25 = io_in_a_bits_address ^ 9'h044;
	wire [9:0] _T_26 = {1'b0, $signed(_T_25)};
	wire [9:0] _T_28 = $signed(_T_26) & -10'sh00c;
	wire _T_29 = $signed(_T_28) == 10'sh000;
	wire [8:0] _T_30 = io_in_a_bits_address ^ 9'h058;
	wire [9:0] _T_31 = {1'b0, $signed(_T_30)};
	wire [9:0] _T_33 = $signed(_T_31) & -10'sh008;
	wire _T_34 = $signed(_T_33) == 10'sh000;
	wire [8:0] _T_35 = io_in_a_bits_address ^ 9'h060;
	wire [9:0] _T_36 = {1'b0, $signed(_T_35)};
	wire [9:0] _T_38 = $signed(_T_36) & -10'sh020;
	wire _T_39 = $signed(_T_38) == 10'sh000;
	wire [8:0] _T_40 = io_in_a_bits_address ^ 9'h080;
	wire [9:0] _T_41 = {1'b0, $signed(_T_40)};
	wire [9:0] _T_43 = $signed(_T_41) & -10'sh080;
	wire _T_44 = $signed(_T_43) == 10'sh000;
	wire [8:0] _T_45 = io_in_a_bits_address ^ 9'h100;
	wire [9:0] _T_46 = {1'b0, $signed(_T_45)};
	wire [9:0] _T_48 = $signed(_T_46) & -10'sh100;
	wire _T_49 = $signed(_T_48) == 10'sh000;
	wire _T_54 = ((((_T_24 | _T_29) | _T_34) | _T_39) | _T_44) | _T_49;
	wire _T_116 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_120 = ~io_in_a_bits_mask;
	wire _T_121 = _T_120 == 4'h0;
	wire _T_125 = ~io_in_a_bits_corrupt;
	wire _T_129 = io_in_a_bits_opcode == 3'h7;
	wire _T_234 = io_in_a_bits_param != 3'h0;
	wire _T_247 = io_in_a_bits_opcode == 3'h4;
	wire _T_248 = 2'h2 == io_in_a_bits_size;
	wire _T_250 = _T_248 & _source_ok_T;
	wire _T_256 = io_in_a_bits_size <= 2'h2;
	wire _T_294 = _T_256 & _T_54;
	wire _T_305 = io_in_a_bits_param == 3'h0;
	wire _T_309 = io_in_a_bits_mask == mask;
	wire _T_317 = io_in_a_bits_opcode == 3'h0;
	wire _T_363 = _T_250 & _T_294;
	wire _T_381 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_440 = ~mask;
	wire [3:0] _T_441 = io_in_a_bits_mask & _T_440;
	wire _T_442 = _T_441 == 4'h0;
	wire _T_446 = io_in_a_bits_opcode == 3'h2;
	wire _T_498 = io_in_a_bits_param <= 3'h4;
	wire _T_506 = io_in_a_bits_opcode == 3'h3;
	wire _T_558 = io_in_a_bits_param <= 3'h3;
	wire _T_566 = io_in_a_bits_opcode == 3'h5;
	wire _T_618 = io_in_a_bits_param <= 3'h1;
	wire _T_630 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_1 = ~io_in_d_bits_source;
	wire _T_634 = io_in_d_bits_opcode == 3'h6;
	wire _T_638 = io_in_d_bits_size >= 2'h2;
	wire _T_654 = io_in_d_bits_opcode == 3'h4;
	wire _T_682 = io_in_d_bits_opcode == 3'h5;
	wire _T_711 = io_in_d_bits_opcode == 3'h0;
	wire _T_728 = io_in_d_bits_opcode == 3'h1;
	wire _T_746 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [1:0] size;
	reg source;
	reg [8:0] address;
	wire _T_776 = io_in_a_valid & ~a_first;
	wire _T_777 = io_in_a_bits_opcode == opcode;
	wire _T_781 = io_in_a_bits_param == param;
	wire _T_785 = io_in_a_bits_size == size;
	wire _T_789 = io_in_a_bits_source == source;
	wire _T_793 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] size_1;
	reg source_1;
	wire _T_800 = io_in_d_valid & ~d_first;
	wire _T_801 = io_in_d_bits_opcode == opcode_1;
	wire _T_809 = io_in_d_bits_size == size_1;
	wire _T_813 = io_in_d_bits_source == source_1;
	reg inflight;
	reg [3:0] inflight_opcodes;
	reg [3:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [3:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [15:0] _GEN_73 = {12'd0, _a_opcode_lookup_T_1};
	wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5;
	wire [15:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[15:1]};
	wire [3:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [15:0] _GEN_76 = {12'd0, _a_size_lookup_T_1};
	wire [15:0] _a_size_lookup_T_6 = _GEN_76 & _a_opcode_lookup_T_5;
	wire [15:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[15:1]};
	wire _T_827 = io_in_a_valid & a_first_1;
	wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source;
	wire _T_830 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1;
	wire [2:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [3:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [18:0] _GEN_1 = {15'd0, a_opcodes_set_interm};
	wire [18:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? _a_sizes_set_interm_T_1 : 3'h0);
	wire [17:0] _GEN_2 = {15'd0, a_sizes_set_interm};
	wire [17:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire _T_834 = ~(inflight >> io_in_a_bits_source);
	wire [1:0] _GEN_16 = (a_first_done & a_first_1 ? _a_set_wo_ready_T : 2'h0);
	wire [18:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 19'h00000);
	wire [17:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 18'h00000);
	wire _T_838 = io_in_d_valid & d_first_1;
	wire _T_840 = ~_T_634;
	wire _T_841 = (io_in_d_valid & d_first_1) & ~_T_634;
	wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source;
	wire [30:0] _GEN_3 = {15'd0, _a_opcode_lookup_T_5};
	wire [30:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [1:0] _GEN_22 = ((d_first_done & d_first_1) & _T_840 ? _d_clr_wo_ready_T : 2'h0);
	wire [30:0] _GEN_23 = ((d_first_done & d_first_1) & _T_840 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_827 & (io_in_a_bits_source == io_in_d_bits_source);
	wire _T_853 = (inflight >> io_in_d_bits_source) | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_858 = io_in_d_bits_opcode == _GEN_40;
	wire _T_859 = (io_in_d_bits_opcode == _GEN_32) | _T_858;
	wire _T_863 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_870 = io_in_d_bits_opcode == _GEN_56;
	wire _T_871 = (io_in_d_bits_opcode == _GEN_48) | _T_870;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {2'd0, io_in_d_bits_size};
	wire _T_875 = _GEN_82 == a_size_lookup;
	wire _T_885 = (((_T_838 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_840;
	wire _T_887 = ~io_in_d_ready | io_in_a_ready;
	wire a_set = _GEN_16[0];
	wire d_clr = _GEN_22[0];
	wire [3:0] a_opcodes_set = _GEN_19[3:0];
	wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [3:0] d_opcodes_clr = _GEN_23[3:0];
	wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [3:0] a_sizes_set = _GEN_20[3:0];
	wire [3:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [3:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_896 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [3:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [3:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [15:0] _GEN_87 = {12'd0, _c_size_lookup_T_1};
	wire [15:0] _c_size_lookup_T_6 = _GEN_87 & _a_opcode_lookup_T_5;
	wire [15:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[15:1]};
	wire _T_922 = (io_in_d_valid & d_first_2) & _T_634;
	wire [30:0] _GEN_68 = ((d_first_done & d_first_2) & _T_634 ? _d_opcodes_clr_T_5 : 31'h00000000);
	wire _T_930 = 1'h0 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_940 = _GEN_82 == c_size_lookup;
	wire [3:0] d_opcodes_clr_1 = _GEN_68[3:0];
	wire [3:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [3:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			param <= io_in_a_bits_param;
		if (a_first_done & a_first)
			size <= io_in_a_bits_size;
		if (a_first_done & a_first)
			source <= io_in_a_bits_source;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 1'h0;
		else
			inflight <= (inflight | a_set) & ~d_clr;
		if (reset)
			inflight_opcodes <= 4'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 4'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_sizes_1 <= 4'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
	end
endmodule
module TLMonitor_42 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [1:0] io_in_a_bits_size;
	input [7:0] io_in_a_bits_source;
	input [11:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_size;
	input [7:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_4 = io_in_a_bits_source <= 8'h9f;
	wire [4:0] _is_aligned_mask_T_1 = 5'h03 << io_in_a_bits_size;
	wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0];
	wire [11:0] _GEN_71 = {10'd0, is_aligned_mask};
	wire [11:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 12'h000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 2'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_10 = ~_source_ok_T_4;
	wire [12:0] _T_12 = {1'b0, $signed(io_in_a_bits_address)};
	wire _T_20 = io_in_a_bits_opcode == 3'h6;
	wire [12:0] _T_36 = $signed(_T_12) & 13'sh1000;
	wire _T_37 = $signed(_T_36) == 13'sh0000;
	wire _T_69 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_73 = ~io_in_a_bits_mask;
	wire _T_74 = _T_73 == 4'h0;
	wire _T_78 = ~io_in_a_bits_corrupt;
	wire _T_82 = io_in_a_bits_opcode == 3'h7;
	wire _T_135 = io_in_a_bits_param != 3'h0;
	wire _T_148 = io_in_a_bits_opcode == 3'h4;
	wire _T_164 = io_in_a_bits_size <= 2'h2;
	wire _T_172 = _T_164 & _T_37;
	wire _T_183 = io_in_a_bits_param == 3'h0;
	wire _T_187 = io_in_a_bits_mask == mask;
	wire _T_195 = io_in_a_bits_opcode == 3'h0;
	wire _T_218 = _source_ok_T_4 & _T_172;
	wire _T_236 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_273 = ~mask;
	wire [3:0] _T_274 = io_in_a_bits_mask & _T_273;
	wire _T_275 = _T_274 == 4'h0;
	wire _T_279 = io_in_a_bits_opcode == 3'h2;
	wire _T_309 = io_in_a_bits_param <= 3'h4;
	wire _T_317 = io_in_a_bits_opcode == 3'h3;
	wire _T_347 = io_in_a_bits_param <= 3'h3;
	wire _T_355 = io_in_a_bits_opcode == 3'h5;
	wire _T_385 = io_in_a_bits_param <= 3'h1;
	wire _T_397 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_10 = io_in_d_bits_source <= 8'h9f;
	wire _T_401 = io_in_d_bits_opcode == 3'h6;
	wire _T_405 = io_in_d_bits_size >= 2'h2;
	wire _T_421 = io_in_d_bits_opcode == 3'h4;
	wire _T_449 = io_in_d_bits_opcode == 3'h5;
	wire _T_478 = io_in_d_bits_opcode == 3'h0;
	wire _T_495 = io_in_d_bits_opcode == 3'h1;
	wire _T_513 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [1:0] size;
	reg [7:0] source;
	reg [11:0] address;
	wire _T_543 = io_in_a_valid & ~a_first;
	wire _T_544 = io_in_a_bits_opcode == opcode;
	wire _T_548 = io_in_a_bits_param == param;
	wire _T_552 = io_in_a_bits_size == size;
	wire _T_556 = io_in_a_bits_source == source;
	wire _T_560 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] size_1;
	reg [7:0] source_1;
	wire _T_567 = io_in_d_valid & ~d_first;
	wire _T_568 = io_in_d_bits_opcode == opcode_1;
	wire _T_576 = io_in_d_bits_size == size_1;
	wire _T_580 = io_in_d_bits_source == source_1;
	reg [159:0] inflight;
	reg [639:0] inflight_opcodes;
	reg [639:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [10:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [639:0] _GEN_73 = {624'd0, _a_opcode_lookup_T_5};
	wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [639:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[639:1]};
	wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [639:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[639:1]};
	wire _T_594 = io_in_a_valid & a_first_1;
	wire [255:0] _a_set_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_a_bits_source;
	wire _T_597 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1;
	wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [10:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [2050:0] _GEN_1 = {2047'd0, a_opcodes_set_interm};
	wire [2050:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? _a_sizes_set_interm_T_1 : 3'h0);
	wire [2049:0] _GEN_2 = {2047'd0, a_sizes_set_interm};
	wire [2049:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [159:0] _T_599 = inflight >> io_in_a_bits_source;
	wire _T_601 = ~_T_599[0];
	wire [255:0] _GEN_16 = (a_first_done & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2050:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 2051'h0);
	wire [2049:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 2050'h0);
	wire _T_605 = io_in_d_valid & d_first_1;
	wire _T_607 = ~_T_401;
	wire _T_608 = (io_in_d_valid & d_first_1) & ~_T_401;
	wire [255:0] _d_clr_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_d_bits_source;
	wire [2062:0] _GEN_3 = {2047'd0, _a_opcode_lookup_T_5};
	wire [2062:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [255:0] _GEN_22 = ((d_first_done & d_first_1) & _T_607 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_23 = ((d_first_done & d_first_1) & _T_607 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_594 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [159:0] _T_618 = inflight >> io_in_d_bits_source;
	wire _T_620 = _T_618[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_625 = io_in_d_bits_opcode == _GEN_40;
	wire _T_626 = (io_in_d_bits_opcode == _GEN_32) | _T_625;
	wire _T_630 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_637 = io_in_d_bits_opcode == _GEN_56;
	wire _T_638 = (io_in_d_bits_opcode == _GEN_48) | _T_637;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {2'd0, io_in_d_bits_size};
	wire _T_642 = _GEN_82 == a_size_lookup;
	wire _T_652 = (((_T_605 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_607;
	wire _T_654 = ~io_in_d_ready | io_in_a_ready;
	wire [159:0] a_set = _GEN_16[159:0];
	wire [159:0] _inflight_T = inflight | a_set;
	wire [159:0] d_clr = _GEN_22[159:0];
	wire [159:0] _inflight_T_1 = ~d_clr;
	wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [639:0] a_opcodes_set = _GEN_19[639:0];
	wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [639:0] d_opcodes_clr = _GEN_23[639:0];
	wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [639:0] a_sizes_set = _GEN_20[639:0];
	wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_663 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [159:0] inflight_1;
	reg [639:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [639:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[639:1]};
	wire _T_689 = (io_in_d_valid & d_first_2) & _T_401;
	wire [255:0] _GEN_67 = ((d_first_done & d_first_2) & _T_401 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_68 = ((d_first_done & d_first_2) & _T_401 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire [159:0] _T_697 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_707 = _GEN_82 == c_size_lookup;
	wire [159:0] d_clr_1 = _GEN_67[159:0];
	wire [159:0] _inflight_T_4 = ~d_clr_1;
	wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0];
	wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_727 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			param <= io_in_a_bits_param;
		if (a_first_done & a_first)
			size <= io_in_a_bits_size;
		if (a_first_done & a_first)
			source <= io_in_a_bits_source;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 160'h0000000000000000000000000000000000000000;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 640'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 640'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 160'h0000000000000000000000000000000000000000;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 640'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (d_first_done)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module TLDebugModuleInner (
	clock,
	reset,
	auto_tl_in_a_ready,
	auto_tl_in_a_valid,
	auto_tl_in_a_bits_opcode,
	auto_tl_in_a_bits_param,
	auto_tl_in_a_bits_size,
	auto_tl_in_a_bits_source,
	auto_tl_in_a_bits_address,
	auto_tl_in_a_bits_mask,
	auto_tl_in_a_bits_data,
	auto_tl_in_a_bits_corrupt,
	auto_tl_in_d_ready,
	auto_tl_in_d_valid,
	auto_tl_in_d_bits_opcode,
	auto_tl_in_d_bits_size,
	auto_tl_in_d_bits_source,
	auto_tl_in_d_bits_data,
	auto_dmi_in_a_ready,
	auto_dmi_in_a_valid,
	auto_dmi_in_a_bits_opcode,
	auto_dmi_in_a_bits_param,
	auto_dmi_in_a_bits_size,
	auto_dmi_in_a_bits_source,
	auto_dmi_in_a_bits_address,
	auto_dmi_in_a_bits_mask,
	auto_dmi_in_a_bits_data,
	auto_dmi_in_a_bits_corrupt,
	auto_dmi_in_d_ready,
	auto_dmi_in_d_valid,
	auto_dmi_in_d_bits_opcode,
	auto_dmi_in_d_bits_size,
	auto_dmi_in_d_bits_source,
	auto_dmi_in_d_bits_data,
	io_dmactive,
	io_innerCtrl_ready,
	io_innerCtrl_valid,
	io_innerCtrl_bits_resumereq,
	io_innerCtrl_bits_hartsel,
	io_innerCtrl_bits_ackhavereset,
	io_innerCtrl_bits_hrmask_0,
	io_hgDebugInt_0,
	io_hartIsInReset_0
);
	input clock;
	input reset;
	output wire auto_tl_in_a_ready;
	input auto_tl_in_a_valid;
	input [2:0] auto_tl_in_a_bits_opcode;
	input [2:0] auto_tl_in_a_bits_param;
	input [1:0] auto_tl_in_a_bits_size;
	input [7:0] auto_tl_in_a_bits_source;
	input [11:0] auto_tl_in_a_bits_address;
	input [3:0] auto_tl_in_a_bits_mask;
	input [31:0] auto_tl_in_a_bits_data;
	input auto_tl_in_a_bits_corrupt;
	input auto_tl_in_d_ready;
	output wire auto_tl_in_d_valid;
	output wire [2:0] auto_tl_in_d_bits_opcode;
	output wire [1:0] auto_tl_in_d_bits_size;
	output wire [7:0] auto_tl_in_d_bits_source;
	output wire [31:0] auto_tl_in_d_bits_data;
	output wire auto_dmi_in_a_ready;
	input auto_dmi_in_a_valid;
	input [2:0] auto_dmi_in_a_bits_opcode;
	input [2:0] auto_dmi_in_a_bits_param;
	input [1:0] auto_dmi_in_a_bits_size;
	input auto_dmi_in_a_bits_source;
	input [8:0] auto_dmi_in_a_bits_address;
	input [3:0] auto_dmi_in_a_bits_mask;
	input [31:0] auto_dmi_in_a_bits_data;
	input auto_dmi_in_a_bits_corrupt;
	input auto_dmi_in_d_ready;
	output wire auto_dmi_in_d_valid;
	output wire [2:0] auto_dmi_in_d_bits_opcode;
	output wire [1:0] auto_dmi_in_d_bits_size;
	output wire auto_dmi_in_d_bits_source;
	output wire [31:0] auto_dmi_in_d_bits_data;
	input io_dmactive;
	output wire io_innerCtrl_ready;
	input io_innerCtrl_valid;
	input io_innerCtrl_bits_resumereq;
	input [9:0] io_innerCtrl_bits_hartsel;
	input io_innerCtrl_bits_ackhavereset;
	input io_innerCtrl_bits_hrmask_0;
	output wire io_hgDebugInt_0;
	input io_hartIsInReset_0;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [1:0] monitor_io_in_a_bits_size;
	wire monitor_io_in_a_bits_source;
	wire [8:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_size;
	wire monitor_io_in_d_bits_source;
	wire monitor_1_clock;
	wire monitor_1_reset;
	wire monitor_1_io_in_a_ready;
	wire monitor_1_io_in_a_valid;
	wire [2:0] monitor_1_io_in_a_bits_opcode;
	wire [2:0] monitor_1_io_in_a_bits_param;
	wire [1:0] monitor_1_io_in_a_bits_size;
	wire [7:0] monitor_1_io_in_a_bits_source;
	wire [11:0] monitor_1_io_in_a_bits_address;
	wire [3:0] monitor_1_io_in_a_bits_mask;
	wire monitor_1_io_in_a_bits_corrupt;
	wire monitor_1_io_in_d_ready;
	wire monitor_1_io_in_d_valid;
	wire [2:0] monitor_1_io_in_d_bits_opcode;
	wire [1:0] monitor_1_io_in_d_bits_size;
	wire [7:0] monitor_1_io_in_d_bits_source;
	wire hartIsInResetSync_0_debug_hartReset_0_clock;
	wire hartIsInResetSync_0_debug_hartReset_0_reset;
	wire hartIsInResetSync_0_debug_hartReset_0_io_d;
	wire hartIsInResetSync_0_debug_hartReset_0_io_q;
	reg haltedBitRegs;
	reg resumeReqRegs;
	reg haveResetBitRegs;
	wire hamaskWrSel_0 = io_innerCtrl_bits_hartsel == 10'h000;
	reg hrmaskReg_0;
	wire _T_1 = ~io_dmactive;
	wire _T_4 = io_innerCtrl_ready & io_innerCtrl_valid;
	reg hrDebugIntReg_0;
	wire _T_10 = ~haltedBitRegs;
	wire _T_11 = hrDebugIntReg_0 & _T_10;
	wire hartIsInResetSync_0 = hartIsInResetSync_0_debug_hartReset_0_io_q;
	wire _T_12 = hartIsInResetSync_0 | _T_11;
	wire _T_13 = hrmaskReg_0 & _T_12;
	wire resumereq = _T_4 & io_innerCtrl_bits_resumereq;
	wire _resumeAcks_T_1 = ~hamaskWrSel_0;
	wire resumeAcks = (resumereq ? ~resumeReqRegs & ~hamaskWrSel_0 : ~resumeReqRegs);
	wire [31:0] haltedStatus_0 = {31'd0, haltedBitRegs};
	wire haltedSummary = |haltedStatus_0;
	wire [31:0] HALTSUM1RdData_haltsum1 = {31'd0, haltedSummary};
	reg [2:0] ABSTRACTCSReg_cmderr;
	wire in_bits_read = auto_dmi_in_a_bits_opcode == 3'h4;
	wire [6:0] in_bits_index = auto_dmi_in_a_bits_address[8:2];
	wire [4:0] out_iindex = {in_bits_index[5], in_bits_index[3], in_bits_index[2], in_bits_index[1], in_bits_index[0]};
	wire [6:0] out_findex = in_bits_index & 7'h50;
	wire _out_T_44 = out_findex == 7'h00;
	wire _out_T_2 = out_findex == 7'h10;
	wire _out_T_20 = out_findex == 7'h40;
	wire [31:0] _out_backSel_T = 32'h00000001 << out_iindex;
	wire out_backSel_6 = _out_backSel_T[6];
	wire out_woready__61 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_6) & (out_findex == 7'h10);
	wire [7:0] _out_backMask_T_11 = (auto_dmi_in_a_bits_mask[3] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_9 = (auto_dmi_in_a_bits_mask[2] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_7 = (auto_dmi_in_a_bits_mask[1] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_5 = (auto_dmi_in_a_bits_mask[0] ? 8'hff : 8'h00);
	wire [31:0] out_backMask = {_out_backMask_T_11, _out_backMask_T_9, _out_backMask_T_7, _out_backMask_T_5};
	wire out_womask_61 = &out_backMask[10:8];
	wire out_f_woready_61 = out_woready__61 & out_womask_61;
	reg [1:0] ctrlStateReg;
	wire ABSTRACTCSWrEnLegal = ctrlStateReg == 2'h0;
	wire ABSTRACTCSWrEn = out_f_woready_61 & ABSTRACTCSWrEnLegal;
	wire [2:0] ABSTRACTCSWrData_cmderr = auto_dmi_in_a_bits_data[10:8];
	wire [2:0] _ABSTRACTCSReg_cmderr_T = ~ABSTRACTCSWrData_cmderr;
	wire [2:0] _ABSTRACTCSReg_cmderr_T_1 = ABSTRACTCSReg_cmderr & _ABSTRACTCSReg_cmderr_T;
	wire [2:0] _GEN_37 = (ABSTRACTCSWrEn ? _ABSTRACTCSReg_cmderr_T_1 : ABSTRACTCSReg_cmderr);
	wire _T_1383 = ctrlStateReg == 2'h1;
	reg [7:0] COMMANDRdData_cmdtype;
	wire commandRegIsAccessRegister = COMMANDRdData_cmdtype == 8'h00;
	reg [23:0] COMMANDRdData_control;
	wire [31:0] _accessRegisterCommandReg_T = {COMMANDRdData_cmdtype, COMMANDRdData_control};
	wire accessRegisterCommandReg_transfer = _accessRegisterCommandReg_T[17];
	wire accessRegisterCommandReg_write = _accessRegisterCommandReg_T[16];
	wire [15:0] accessRegisterCommandReg_regno = _accessRegisterCommandReg_T[15:0];
	wire [2:0] accessRegisterCommandReg_size = _accessRegisterCommandReg_T[22:20];
	wire accessRegIsLegalSize = (accessRegisterCommandReg_size == 3'h2) | (accessRegisterCommandReg_size == 3'h3);
	wire accessRegIsGPR = ((accessRegisterCommandReg_regno >= 16'h1000) & (accessRegisterCommandReg_regno <= 16'h101f)) & accessRegIsLegalSize;
	wire _GEN_3614 = (~accessRegisterCommandReg_transfer | accessRegIsGPR ? 1'h0 : 1'h1);
	wire commandRegIsUnsupported = (commandRegIsAccessRegister ? _GEN_3614 : 1'h1);
	wire _GEN_3615 = (~accessRegisterCommandReg_transfer | accessRegIsGPR) & _T_10;
	wire commandRegBadHaltResume = commandRegIsAccessRegister & _GEN_3615;
	wire _GEN_3631 = (commandRegIsUnsupported ? 1'h0 : commandRegBadHaltResume);
	wire _GEN_3644 = (ctrlStateReg == 2'h1) & _GEN_3631;
	wire errorHaltResume = (ABSTRACTCSWrEnLegal ? 1'h0 : _GEN_3644);
	wire [2:0] _GEN_38 = (errorHaltResume ? 3'h4 : _GEN_37);
	wire out_backSel_7 = _out_backSel_T[7];
	wire out_woready__86 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_7) & (out_findex == 7'h10);
	wire out_womask_86 = &out_backMask;
	wire out_f_woready_86 = out_woready__86 & out_womask_86;
	wire COMMANDWrEn = out_f_woready_86 & ABSTRACTCSWrEnLegal;
	wire [31:0] COMMANDWrDataVal = (out_f_woready_86 ? auto_dmi_in_a_bits_data : 32'h00000000);
	wire [7:0] COMMANDWrData_cmdtype = COMMANDWrDataVal[31:24];
	wire commandWrIsAccessRegister = COMMANDWrData_cmdtype == 8'h00;
	wire _wrAccessRegisterCommand_T_1 = ABSTRACTCSReg_cmderr == 3'h0;
	wire wrAccessRegisterCommand = (COMMANDWrEn & commandWrIsAccessRegister) & (ABSTRACTCSReg_cmderr == 3'h0);
	wire out_backSel_4 = _out_backSel_T[4];
	wire out_woready__92 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_4) & (out_findex == 7'h00);
	wire out_womask_92 = &out_backMask[7:0];
	wire out_f_woready_92 = out_woready__92 & out_womask_92;
	wire out_roready__92 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_4) & (out_findex == 7'h00);
	wire out_romask_92 = |out_backMask[7:0];
	wire out_f_roready_92 = out_roready__92 & out_romask_92;
	wire dmiAbstractDataAccessVec_0 = out_f_woready_92 | out_f_roready_92;
	reg [11:0] ABSTRACTAUTOReg_autoexecdata;
	wire autoexecData_0 = dmiAbstractDataAccessVec_0 & ABSTRACTAUTOReg_autoexecdata[0];
	wire out_backSel_16 = _out_backSel_T[16];
	wire out_woready__27 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_16) & (out_findex == 7'h00);
	wire out_f_woready_27 = out_woready__27 & out_womask_92;
	wire out_roready__27 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_16) & (out_findex == 7'h00);
	wire out_f_roready_27 = out_roready__27 & out_romask_92;
	wire dmiProgramBufferAccessVec_0 = out_f_woready_27 | out_f_roready_27;
	reg [15:0] ABSTRACTAUTOReg_autoexecprogbuf;
	wire autoexecProg_0 = dmiProgramBufferAccessVec_0 & ABSTRACTAUTOReg_autoexecprogbuf[0];
	wire out_backSel_17 = _out_backSel_T[17];
	wire out_woready__19 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_17) & (out_findex == 7'h00);
	wire out_f_woready_19 = out_woready__19 & out_womask_92;
	wire out_roready__19 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_17) & (out_findex == 7'h00);
	wire out_f_roready_19 = out_roready__19 & out_romask_92;
	wire dmiProgramBufferAccessVec_4 = out_f_woready_19 | out_f_roready_19;
	wire autoexecProg_1 = dmiProgramBufferAccessVec_4 & ABSTRACTAUTOReg_autoexecprogbuf[1];
	wire out_backSel_18 = _out_backSel_T[18];
	wire out_woready__31 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_18) & (out_findex == 7'h00);
	wire out_f_woready_31 = out_woready__31 & out_womask_92;
	wire out_roready__31 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_18) & (out_findex == 7'h00);
	wire out_f_roready_31 = out_roready__31 & out_romask_92;
	wire dmiProgramBufferAccessVec_8 = out_f_woready_31 | out_f_roready_31;
	wire autoexecProg_2 = dmiProgramBufferAccessVec_8 & ABSTRACTAUTOReg_autoexecprogbuf[2];
	wire out_backSel_19 = _out_backSel_T[19];
	wire out_woready__74 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_19) & (out_findex == 7'h00);
	wire out_f_woready_74 = out_woready__74 & out_womask_92;
	wire out_roready__74 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_19) & (out_findex == 7'h00);
	wire out_f_roready_74 = out_roready__74 & out_romask_92;
	wire dmiProgramBufferAccessVec_12 = out_f_woready_74 | out_f_roready_74;
	wire autoexecProg_3 = dmiProgramBufferAccessVec_12 & ABSTRACTAUTOReg_autoexecprogbuf[3];
	wire out_backSel_20 = _out_backSel_T[20];
	wire out_woready__87 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_20) & (out_findex == 7'h00);
	wire out_f_woready_87 = out_woready__87 & out_womask_92;
	wire out_roready__87 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_20) & (out_findex == 7'h00);
	wire out_f_roready_87 = out_roready__87 & out_romask_92;
	wire dmiProgramBufferAccessVec_16 = out_f_woready_87 | out_f_roready_87;
	wire autoexecProg_4 = dmiProgramBufferAccessVec_16 & ABSTRACTAUTOReg_autoexecprogbuf[4];
	wire out_backSel_21 = _out_backSel_T[21];
	wire out_woready__7 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_21) & (out_findex == 7'h00);
	wire out_f_woready_7 = out_woready__7 & out_womask_92;
	wire out_roready__7 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_21) & (out_findex == 7'h00);
	wire out_f_roready_7 = out_roready__7 & out_romask_92;
	wire dmiProgramBufferAccessVec_20 = out_f_woready_7 | out_f_roready_7;
	wire autoexecProg_5 = dmiProgramBufferAccessVec_20 & ABSTRACTAUTOReg_autoexecprogbuf[5];
	wire out_backSel_22 = _out_backSel_T[22];
	wire out_woready__15 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_22) & (out_findex == 7'h00);
	wire out_f_woready_15 = out_woready__15 & out_womask_92;
	wire out_roready__15 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_22) & (out_findex == 7'h00);
	wire out_f_roready_15 = out_roready__15 & out_romask_92;
	wire dmiProgramBufferAccessVec_24 = out_f_woready_15 | out_f_roready_15;
	wire autoexecProg_6 = dmiProgramBufferAccessVec_24 & ABSTRACTAUTOReg_autoexecprogbuf[6];
	wire out_backSel_23 = _out_backSel_T[23];
	wire out_woready__70 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_23) & (out_findex == 7'h00);
	wire out_f_woready_70 = out_woready__70 & out_womask_92;
	wire out_roready__70 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_23) & (out_findex == 7'h00);
	wire out_f_roready_70 = out_roready__70 & out_romask_92;
	wire dmiProgramBufferAccessVec_28 = out_f_woready_70 | out_f_roready_70;
	wire autoexecProg_7 = dmiProgramBufferAccessVec_28 & ABSTRACTAUTOReg_autoexecprogbuf[7];
	wire out_backSel_24 = _out_backSel_T[24];
	wire out_woready__82 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_24) & (out_findex == 7'h00);
	wire out_f_woready_82 = out_woready__82 & out_womask_92;
	wire out_roready__82 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_24) & (out_findex == 7'h00);
	wire out_f_roready_82 = out_roready__82 & out_romask_92;
	wire dmiProgramBufferAccessVec_32 = out_f_woready_82 | out_f_roready_82;
	wire autoexecProg_8 = dmiProgramBufferAccessVec_32 & ABSTRACTAUTOReg_autoexecprogbuf[8];
	wire out_backSel_25 = _out_backSel_T[25];
	wire out_woready__23 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_25) & (out_findex == 7'h00);
	wire out_f_woready_23 = out_woready__23 & out_womask_92;
	wire out_roready__23 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_25) & (out_findex == 7'h00);
	wire out_f_roready_23 = out_roready__23 & out_romask_92;
	wire dmiProgramBufferAccessVec_36 = out_f_woready_23 | out_f_roready_23;
	wire autoexecProg_9 = dmiProgramBufferAccessVec_36 & ABSTRACTAUTOReg_autoexecprogbuf[9];
	wire out_backSel_26 = _out_backSel_T[26];
	wire out_woready__0 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_26) & (out_findex == 7'h00);
	wire out_f_woready = out_woready__0 & out_womask_92;
	wire out_roready__0 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_26) & (out_findex == 7'h00);
	wire out_f_roready = out_roready__0 & out_romask_92;
	wire dmiProgramBufferAccessVec_40 = out_f_woready | out_f_roready;
	wire autoexecProg_10 = dmiProgramBufferAccessVec_40 & ABSTRACTAUTOReg_autoexecprogbuf[10];
	wire out_backSel_27 = _out_backSel_T[27];
	wire out_woready__78 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_27) & (out_findex == 7'h00);
	wire out_f_woready_78 = out_woready__78 & out_womask_92;
	wire out_roready__78 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_27) & (out_findex == 7'h00);
	wire out_f_roready_78 = out_roready__78 & out_romask_92;
	wire dmiProgramBufferAccessVec_44 = out_f_woready_78 | out_f_roready_78;
	wire autoexecProg_11 = dmiProgramBufferAccessVec_44 & ABSTRACTAUTOReg_autoexecprogbuf[11];
	wire out_backSel_28 = _out_backSel_T[28];
	wire out_woready__66 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_28) & (out_findex == 7'h00);
	wire out_f_woready_66 = out_woready__66 & out_womask_92;
	wire out_roready__66 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_28) & (out_findex == 7'h00);
	wire out_f_roready_66 = out_roready__66 & out_romask_92;
	wire dmiProgramBufferAccessVec_48 = out_f_woready_66 | out_f_roready_66;
	wire autoexecProg_12 = dmiProgramBufferAccessVec_48 & ABSTRACTAUTOReg_autoexecprogbuf[12];
	wire out_backSel_29 = _out_backSel_T[29];
	wire out_woready__35 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_29) & (out_findex == 7'h00);
	wire out_f_woready_35 = out_woready__35 & out_womask_92;
	wire out_roready__35 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_29) & (out_findex == 7'h00);
	wire out_f_roready_35 = out_roready__35 & out_romask_92;
	wire dmiProgramBufferAccessVec_52 = out_f_woready_35 | out_f_roready_35;
	wire autoexecProg_13 = dmiProgramBufferAccessVec_52 & ABSTRACTAUTOReg_autoexecprogbuf[13];
	wire out_backSel_30 = _out_backSel_T[30];
	wire out_woready__11 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_30) & (out_findex == 7'h00);
	wire out_f_woready_11 = out_woready__11 & out_womask_92;
	wire out_roready__11 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_30) & (out_findex == 7'h00);
	wire out_f_roready_11 = out_roready__11 & out_romask_92;
	wire dmiProgramBufferAccessVec_56 = out_f_woready_11 | out_f_roready_11;
	wire autoexecProg_14 = dmiProgramBufferAccessVec_56 & ABSTRACTAUTOReg_autoexecprogbuf[14];
	wire out_backSel_31 = _out_backSel_T[31];
	wire out_woready__96 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_31) & (out_findex == 7'h00);
	wire out_f_woready_96 = out_woready__96 & out_womask_92;
	wire out_roready__96 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & in_bits_read) & out_backSel_31) & (out_findex == 7'h00);
	wire out_f_roready_96 = out_roready__96 & out_romask_92;
	wire dmiProgramBufferAccessVec_60 = out_f_woready_96 | out_f_roready_96;
	wire autoexecProg_15 = dmiProgramBufferAccessVec_60 & ABSTRACTAUTOReg_autoexecprogbuf[15];
	wire autoexec = autoexecData_0 | (((((((((((((((autoexecProg_0 | autoexecProg_1) | autoexecProg_2) | autoexecProg_3) | autoexecProg_4) | autoexecProg_5) | autoexecProg_6) | autoexecProg_7) | autoexecProg_8) | autoexecProg_9) | autoexecProg_10) | autoexecProg_11) | autoexecProg_12) | autoexecProg_13) | autoexecProg_14) | autoexecProg_15);
	wire regAccessRegisterCommand = (autoexec & commandRegIsAccessRegister) & _wrAccessRegisterCommand_T_1;
	wire commandWrIsUnsupported = COMMANDWrEn & ~commandWrIsAccessRegister;
	wire _T_1382 = autoexec & commandRegIsUnsupported;
	wire _GEN_3621 = commandWrIsUnsupported | _T_1382;
	wire _GEN_3623 = (wrAccessRegisterCommand | regAccessRegisterCommand ? 1'h0 : _GEN_3621);
	wire _GEN_3642 = (ctrlStateReg == 2'h1) & commandRegIsUnsupported;
	wire errorUnsupported = (ABSTRACTCSWrEnLegal ? _GEN_3623 : _GEN_3642);
	wire _T_1384 = ctrlStateReg == 2'h2;
	wire in_1_bits_read = auto_tl_in_a_bits_opcode == 3'h4;
	wire [9:0] in_1_bits_index = auto_tl_in_a_bits_address[11:2];
	wire [8:0] out_iindex_1 = {in_1_bits_index[8], in_1_bits_index[7], in_1_bits_index[6], in_1_bits_index[5], in_1_bits_index[4], in_1_bits_index[3], in_1_bits_index[2], in_1_bits_index[1], in_1_bits_index[0]};
	wire [9:0] out_findex_1 = in_1_bits_index & 10'h200;
	wire _out_T_1122 = out_findex_1 == 10'h000;
	wire _out_T_1642 = out_findex_1 == 10'h200;
	wire [511:0] _out_backSel_T_1 = 512'h1 << out_iindex_1;
	wire out_backSel_67 = _out_backSel_T_1[67];
	wire out_woready_1_841 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_backSel_67) & (out_findex_1 == 10'h000);
	wire [7:0] _out_backMask_T_23 = (auto_tl_in_a_bits_mask[3] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_21 = (auto_tl_in_a_bits_mask[2] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_19 = (auto_tl_in_a_bits_mask[1] ? 8'hff : 8'h00);
	wire [7:0] _out_backMask_T_17 = (auto_tl_in_a_bits_mask[0] ? 8'hff : 8'h00);
	wire [31:0] out_backMask_1 = {_out_backMask_T_23, _out_backMask_T_21, _out_backMask_T_19, _out_backMask_T_17};
	wire out_womask_941 = &out_backMask_1[9:0];
	wire out_f_woready_941 = out_woready_1_841 & out_womask_941;
	wire _GEN_3640 = (ctrlStateReg == 2'h2) & out_f_woready_941;
	wire _GEN_3646 = (ctrlStateReg == 2'h1 ? 1'h0 : _GEN_3640);
	wire errorException = (ABSTRACTCSWrEnLegal ? 1'h0 : _GEN_3646);
	wire _errorBusy_T = ~ABSTRACTCSWrEnLegal;
	wire out_backSel_8 = _out_backSel_T[8];
	wire out_woready__4 = (((auto_dmi_in_a_valid & auto_dmi_in_d_ready) & ~in_bits_read) & out_backSel_8) & (out_findex == 7'h10);
	wire out_womask_4 = &out_backMask[0];
	wire out_f_woready_4 = out_woready__4 & out_womask_4;
	wire _errorBusy_T_3 = out_f_woready_4 & _errorBusy_T;
	wire _errorBusy_T_4 = (out_f_woready_61 & ~ABSTRACTCSWrEnLegal) | _errorBusy_T_3;
	wire out_womask_6 = &out_backMask[31:16];
	wire out_f_woready_6 = out_woready__4 & out_womask_6;
	wire _errorBusy_T_6 = out_f_woready_6 & _errorBusy_T;
	wire _errorBusy_T_7 = _errorBusy_T_4 | _errorBusy_T_6;
	wire _errorBusy_T_9 = out_f_woready_86 & _errorBusy_T;
	wire _errorBusy_T_10 = _errorBusy_T_7 | _errorBusy_T_9;
	wire out_womask_93 = &out_backMask[15:8];
	wire out_f_woready_93 = out_woready__92 & out_womask_93;
	wire out_romask_93 = |out_backMask[15:8];
	wire out_f_roready_93 = out_roready__92 & out_romask_93;
	wire dmiAbstractDataAccessVec_1 = out_f_woready_93 | out_f_roready_93;
	wire out_womask_94 = &out_backMask[23:16];
	wire out_f_woready_94 = out_woready__92 & out_womask_94;
	wire out_romask_94 = |out_backMask[23:16];
	wire out_f_roready_94 = out_roready__92 & out_romask_94;
	wire dmiAbstractDataAccessVec_2 = out_f_woready_94 | out_f_roready_94;
	wire out_womask_95 = &out_backMask[31:24];
	wire out_f_woready_95 = out_woready__92 & out_womask_95;
	wire out_romask_95 = |out_backMask[31:24];
	wire out_f_roready_95 = out_roready__92 & out_romask_95;
	wire dmiAbstractDataAccessVec_3 = out_f_woready_95 | out_f_roready_95;
	wire dmiAbstractDataAccess = ((dmiAbstractDataAccessVec_0 | dmiAbstractDataAccessVec_1) | dmiAbstractDataAccessVec_2) | dmiAbstractDataAccessVec_3;
	wire _errorBusy_T_12 = dmiAbstractDataAccess & _errorBusy_T;
	wire _errorBusy_T_13 = _errorBusy_T_10 | _errorBusy_T_12;
	wire out_f_woready_28 = out_woready__27 & out_womask_93;
	wire out_f_roready_28 = out_roready__27 & out_romask_93;
	wire dmiProgramBufferAccessVec_1 = out_f_woready_28 | out_f_roready_28;
	wire out_f_woready_29 = out_woready__27 & out_womask_94;
	wire out_f_roready_29 = out_roready__27 & out_romask_94;
	wire dmiProgramBufferAccessVec_2 = out_f_woready_29 | out_f_roready_29;
	wire out_f_woready_30 = out_woready__27 & out_womask_95;
	wire out_f_roready_30 = out_roready__27 & out_romask_95;
	wire dmiProgramBufferAccessVec_3 = out_f_woready_30 | out_f_roready_30;
	wire out_f_woready_20 = out_woready__19 & out_womask_93;
	wire out_f_roready_20 = out_roready__19 & out_romask_93;
	wire dmiProgramBufferAccessVec_5 = out_f_woready_20 | out_f_roready_20;
	wire out_f_woready_21 = out_woready__19 & out_womask_94;
	wire out_f_roready_21 = out_roready__19 & out_romask_94;
	wire dmiProgramBufferAccessVec_6 = out_f_woready_21 | out_f_roready_21;
	wire out_f_woready_22 = out_woready__19 & out_womask_95;
	wire out_f_roready_22 = out_roready__19 & out_romask_95;
	wire dmiProgramBufferAccessVec_7 = out_f_woready_22 | out_f_roready_22;
	wire out_f_woready_32 = out_woready__31 & out_womask_93;
	wire out_f_roready_32 = out_roready__31 & out_romask_93;
	wire dmiProgramBufferAccessVec_9 = out_f_woready_32 | out_f_roready_32;
	wire out_f_woready_33 = out_woready__31 & out_womask_94;
	wire out_f_roready_33 = out_roready__31 & out_romask_94;
	wire dmiProgramBufferAccessVec_10 = out_f_woready_33 | out_f_roready_33;
	wire out_f_woready_34 = out_woready__31 & out_womask_95;
	wire out_f_roready_34 = out_roready__31 & out_romask_95;
	wire dmiProgramBufferAccessVec_11 = out_f_woready_34 | out_f_roready_34;
	wire out_f_woready_75 = out_woready__74 & out_womask_93;
	wire out_f_roready_75 = out_roready__74 & out_romask_93;
	wire dmiProgramBufferAccessVec_13 = out_f_woready_75 | out_f_roready_75;
	wire out_f_woready_76 = out_woready__74 & out_womask_94;
	wire out_f_roready_76 = out_roready__74 & out_romask_94;
	wire dmiProgramBufferAccessVec_14 = out_f_woready_76 | out_f_roready_76;
	wire out_f_woready_77 = out_woready__74 & out_womask_95;
	wire out_f_roready_77 = out_roready__74 & out_romask_95;
	wire dmiProgramBufferAccessVec_15 = out_f_woready_77 | out_f_roready_77;
	wire out_f_woready_88 = out_woready__87 & out_womask_93;
	wire out_f_roready_88 = out_roready__87 & out_romask_93;
	wire dmiProgramBufferAccessVec_17 = out_f_woready_88 | out_f_roready_88;
	wire out_f_woready_89 = out_woready__87 & out_womask_94;
	wire out_f_roready_89 = out_roready__87 & out_romask_94;
	wire dmiProgramBufferAccessVec_18 = out_f_woready_89 | out_f_roready_89;
	wire out_f_woready_90 = out_woready__87 & out_womask_95;
	wire out_f_roready_90 = out_roready__87 & out_romask_95;
	wire dmiProgramBufferAccessVec_19 = out_f_woready_90 | out_f_roready_90;
	wire out_f_woready_8 = out_woready__7 & out_womask_93;
	wire out_f_roready_8 = out_roready__7 & out_romask_93;
	wire dmiProgramBufferAccessVec_21 = out_f_woready_8 | out_f_roready_8;
	wire out_f_woready_9 = out_woready__7 & out_womask_94;
	wire out_f_roready_9 = out_roready__7 & out_romask_94;
	wire dmiProgramBufferAccessVec_22 = out_f_woready_9 | out_f_roready_9;
	wire out_f_woready_10 = out_woready__7 & out_womask_95;
	wire out_f_roready_10 = out_roready__7 & out_romask_95;
	wire dmiProgramBufferAccessVec_23 = out_f_woready_10 | out_f_roready_10;
	wire out_f_woready_16 = out_woready__15 & out_womask_93;
	wire out_f_roready_16 = out_roready__15 & out_romask_93;
	wire dmiProgramBufferAccessVec_25 = out_f_woready_16 | out_f_roready_16;
	wire out_f_woready_17 = out_woready__15 & out_womask_94;
	wire out_f_roready_17 = out_roready__15 & out_romask_94;
	wire dmiProgramBufferAccessVec_26 = out_f_woready_17 | out_f_roready_17;
	wire out_f_woready_18 = out_woready__15 & out_womask_95;
	wire out_f_roready_18 = out_roready__15 & out_romask_95;
	wire dmiProgramBufferAccessVec_27 = out_f_woready_18 | out_f_roready_18;
	wire out_f_woready_71 = out_woready__70 & out_womask_93;
	wire out_f_roready_71 = out_roready__70 & out_romask_93;
	wire dmiProgramBufferAccessVec_29 = out_f_woready_71 | out_f_roready_71;
	wire out_f_woready_72 = out_woready__70 & out_womask_94;
	wire out_f_roready_72 = out_roready__70 & out_romask_94;
	wire dmiProgramBufferAccessVec_30 = out_f_woready_72 | out_f_roready_72;
	wire _dmiProgramBufferAccess_T_29 = (((((((((((((((((((((((((((((dmiProgramBufferAccessVec_0 | dmiProgramBufferAccessVec_1) | dmiProgramBufferAccessVec_2) | dmiProgramBufferAccessVec_3) | dmiProgramBufferAccessVec_4) | dmiProgramBufferAccessVec_5) | dmiProgramBufferAccessVec_6) | dmiProgramBufferAccessVec_7) | dmiProgramBufferAccessVec_8) | dmiProgramBufferAccessVec_9) | dmiProgramBufferAccessVec_10) | dmiProgramBufferAccessVec_11) | dmiProgramBufferAccessVec_12) | dmiProgramBufferAccessVec_13) | dmiProgramBufferAccessVec_14) | dmiProgramBufferAccessVec_15) | dmiProgramBufferAccessVec_16) | dmiProgramBufferAccessVec_17) | dmiProgramBufferAccessVec_18) | dmiProgramBufferAccessVec_19) | dmiProgramBufferAccessVec_20) | dmiProgramBufferAccessVec_21) | dmiProgramBufferAccessVec_22) | dmiProgramBufferAccessVec_23) | dmiProgramBufferAccessVec_24) | dmiProgramBufferAccessVec_25) | dmiProgramBufferAccessVec_26) | dmiProgramBufferAccessVec_27) | dmiProgramBufferAccessVec_28) | dmiProgramBufferAccessVec_29) | dmiProgramBufferAccessVec_30;
	wire out_f_woready_73 = out_woready__70 & out_womask_95;
	wire out_f_roready_73 = out_roready__70 & out_romask_95;
	wire dmiProgramBufferAccessVec_31 = out_f_woready_73 | out_f_roready_73;
	wire out_f_woready_83 = out_woready__82 & out_womask_93;
	wire out_f_roready_83 = out_roready__82 & out_romask_93;
	wire dmiProgramBufferAccessVec_33 = out_f_woready_83 | out_f_roready_83;
	wire out_f_woready_84 = out_woready__82 & out_womask_94;
	wire out_f_roready_84 = out_roready__82 & out_romask_94;
	wire dmiProgramBufferAccessVec_34 = out_f_woready_84 | out_f_roready_84;
	wire out_f_woready_85 = out_woready__82 & out_womask_95;
	wire out_f_roready_85 = out_roready__82 & out_romask_95;
	wire dmiProgramBufferAccessVec_35 = out_f_woready_85 | out_f_roready_85;
	wire out_f_woready_24 = out_woready__23 & out_womask_93;
	wire out_f_roready_24 = out_roready__23 & out_romask_93;
	wire dmiProgramBufferAccessVec_37 = out_f_woready_24 | out_f_roready_24;
	wire out_f_woready_25 = out_woready__23 & out_womask_94;
	wire out_f_roready_25 = out_roready__23 & out_romask_94;
	wire dmiProgramBufferAccessVec_38 = out_f_woready_25 | out_f_roready_25;
	wire out_f_woready_26 = out_woready__23 & out_womask_95;
	wire out_f_roready_26 = out_roready__23 & out_romask_95;
	wire dmiProgramBufferAccessVec_39 = out_f_woready_26 | out_f_roready_26;
	wire out_f_woready_1 = out_woready__0 & out_womask_93;
	wire out_f_roready_1 = out_roready__0 & out_romask_93;
	wire dmiProgramBufferAccessVec_41 = out_f_woready_1 | out_f_roready_1;
	wire out_f_woready_2 = out_woready__0 & out_womask_94;
	wire out_f_roready_2 = out_roready__0 & out_romask_94;
	wire dmiProgramBufferAccessVec_42 = out_f_woready_2 | out_f_roready_2;
	wire out_f_woready_3 = out_woready__0 & out_womask_95;
	wire out_f_roready_3 = out_roready__0 & out_romask_95;
	wire dmiProgramBufferAccessVec_43 = out_f_woready_3 | out_f_roready_3;
	wire out_f_woready_79 = out_woready__78 & out_womask_93;
	wire out_f_roready_79 = out_roready__78 & out_romask_93;
	wire dmiProgramBufferAccessVec_45 = out_f_woready_79 | out_f_roready_79;
	wire out_f_woready_80 = out_woready__78 & out_womask_94;
	wire out_f_roready_80 = out_roready__78 & out_romask_94;
	wire dmiProgramBufferAccessVec_46 = out_f_woready_80 | out_f_roready_80;
	wire out_f_woready_81 = out_woready__78 & out_womask_95;
	wire out_f_roready_81 = out_roready__78 & out_romask_95;
	wire dmiProgramBufferAccessVec_47 = out_f_woready_81 | out_f_roready_81;
	wire out_f_woready_67 = out_woready__66 & out_womask_93;
	wire out_f_roready_67 = out_roready__66 & out_romask_93;
	wire dmiProgramBufferAccessVec_49 = out_f_woready_67 | out_f_roready_67;
	wire out_f_woready_68 = out_woready__66 & out_womask_94;
	wire out_f_roready_68 = out_roready__66 & out_romask_94;
	wire dmiProgramBufferAccessVec_50 = out_f_woready_68 | out_f_roready_68;
	wire out_f_woready_69 = out_woready__66 & out_womask_95;
	wire out_f_roready_69 = out_roready__66 & out_romask_95;
	wire dmiProgramBufferAccessVec_51 = out_f_woready_69 | out_f_roready_69;
	wire out_f_woready_36 = out_woready__35 & out_womask_93;
	wire out_f_roready_36 = out_roready__35 & out_romask_93;
	wire dmiProgramBufferAccessVec_53 = out_f_woready_36 | out_f_roready_36;
	wire out_f_woready_37 = out_woready__35 & out_womask_94;
	wire out_f_roready_37 = out_roready__35 & out_romask_94;
	wire dmiProgramBufferAccessVec_54 = out_f_woready_37 | out_f_roready_37;
	wire out_f_woready_38 = out_woready__35 & out_womask_95;
	wire out_f_roready_38 = out_roready__35 & out_romask_95;
	wire dmiProgramBufferAccessVec_55 = out_f_woready_38 | out_f_roready_38;
	wire out_f_woready_12 = out_woready__11 & out_womask_93;
	wire out_f_roready_12 = out_roready__11 & out_romask_93;
	wire dmiProgramBufferAccessVec_57 = out_f_woready_12 | out_f_roready_12;
	wire out_f_woready_13 = out_woready__11 & out_womask_94;
	wire out_f_roready_13 = out_roready__11 & out_romask_94;
	wire dmiProgramBufferAccessVec_58 = out_f_woready_13 | out_f_roready_13;
	wire out_f_woready_14 = out_woready__11 & out_womask_95;
	wire out_f_roready_14 = out_roready__11 & out_romask_95;
	wire dmiProgramBufferAccessVec_59 = out_f_woready_14 | out_f_roready_14;
	wire _dmiProgramBufferAccess_T_59 = (((((((((((((((((((((((((((((_dmiProgramBufferAccess_T_29 | dmiProgramBufferAccessVec_31) | dmiProgramBufferAccessVec_32) | dmiProgramBufferAccessVec_33) | dmiProgramBufferAccessVec_34) | dmiProgramBufferAccessVec_35) | dmiProgramBufferAccessVec_36) | dmiProgramBufferAccessVec_37) | dmiProgramBufferAccessVec_38) | dmiProgramBufferAccessVec_39) | dmiProgramBufferAccessVec_40) | dmiProgramBufferAccessVec_41) | dmiProgramBufferAccessVec_42) | dmiProgramBufferAccessVec_43) | dmiProgramBufferAccessVec_44) | dmiProgramBufferAccessVec_45) | dmiProgramBufferAccessVec_46) | dmiProgramBufferAccessVec_47) | dmiProgramBufferAccessVec_48) | dmiProgramBufferAccessVec_49) | dmiProgramBufferAccessVec_50) | dmiProgramBufferAccessVec_51) | dmiProgramBufferAccessVec_52) | dmiProgramBufferAccessVec_53) | dmiProgramBufferAccessVec_54) | dmiProgramBufferAccessVec_55) | dmiProgramBufferAccessVec_56) | dmiProgramBufferAccessVec_57) | dmiProgramBufferAccessVec_58) | dmiProgramBufferAccessVec_59) | dmiProgramBufferAccessVec_60;
	wire out_f_woready_97 = out_woready__96 & out_womask_93;
	wire out_f_roready_97 = out_roready__96 & out_romask_93;
	wire dmiProgramBufferAccessVec_61 = out_f_woready_97 | out_f_roready_97;
	wire out_f_woready_98 = out_woready__96 & out_womask_94;
	wire out_f_roready_98 = out_roready__96 & out_romask_94;
	wire dmiProgramBufferAccessVec_62 = out_f_woready_98 | out_f_roready_98;
	wire out_f_woready_99 = out_woready__96 & out_womask_95;
	wire out_f_roready_99 = out_roready__96 & out_romask_95;
	wire dmiProgramBufferAccessVec_63 = out_f_woready_99 | out_f_roready_99;
	wire dmiProgramBufferAccess = ((_dmiProgramBufferAccess_T_59 | dmiProgramBufferAccessVec_61) | dmiProgramBufferAccessVec_62) | dmiProgramBufferAccessVec_63;
	wire _errorBusy_T_15 = dmiProgramBufferAccess & _errorBusy_T;
	wire errorBusy = _errorBusy_T_13 | _errorBusy_T_15;
	wire [15:0] ABSTRACTAUTOWrData_autoexecprogbuf = auto_dmi_in_a_bits_data[31:16];
	wire [11:0] ABSTRACTAUTOWrData_autoexecdata = {11'd0, auto_dmi_in_a_bits_data[0]};
	wire [11:0] _ABSTRACTAUTOReg_autoexecdata_T = ABSTRACTAUTOWrData_autoexecdata & 12'h001;
	wire [23:0] COMMANDWrData_control = COMMANDWrDataVal[23:0];
	reg [7:0] abstractDataMem_0;
	reg [7:0] abstractDataMem_1;
	reg [7:0] abstractDataMem_2;
	reg [7:0] abstractDataMem_3;
	reg [7:0] programBufferMem_0;
	reg [7:0] programBufferMem_1;
	reg [7:0] programBufferMem_2;
	reg [7:0] programBufferMem_3;
	reg [7:0] programBufferMem_4;
	reg [7:0] programBufferMem_5;
	reg [7:0] programBufferMem_6;
	reg [7:0] programBufferMem_7;
	reg [7:0] programBufferMem_8;
	reg [7:0] programBufferMem_9;
	reg [7:0] programBufferMem_10;
	reg [7:0] programBufferMem_11;
	reg [7:0] programBufferMem_12;
	reg [7:0] programBufferMem_13;
	reg [7:0] programBufferMem_14;
	reg [7:0] programBufferMem_15;
	reg [7:0] programBufferMem_16;
	reg [7:0] programBufferMem_17;
	reg [7:0] programBufferMem_18;
	reg [7:0] programBufferMem_19;
	reg [7:0] programBufferMem_20;
	reg [7:0] programBufferMem_21;
	reg [7:0] programBufferMem_22;
	reg [7:0] programBufferMem_23;
	reg [7:0] programBufferMem_24;
	reg [7:0] programBufferMem_25;
	reg [7:0] programBufferMem_26;
	reg [7:0] programBufferMem_27;
	reg [7:0] programBufferMem_28;
	reg [7:0] programBufferMem_29;
	reg [7:0] programBufferMem_30;
	reg [7:0] programBufferMem_31;
	reg [7:0] programBufferMem_32;
	reg [7:0] programBufferMem_33;
	reg [7:0] programBufferMem_34;
	reg [7:0] programBufferMem_35;
	reg [7:0] programBufferMem_36;
	reg [7:0] programBufferMem_37;
	reg [7:0] programBufferMem_38;
	reg [7:0] programBufferMem_39;
	reg [7:0] programBufferMem_40;
	reg [7:0] programBufferMem_41;
	reg [7:0] programBufferMem_42;
	reg [7:0] programBufferMem_43;
	reg [7:0] programBufferMem_44;
	reg [7:0] programBufferMem_45;
	reg [7:0] programBufferMem_46;
	reg [7:0] programBufferMem_47;
	reg [7:0] programBufferMem_48;
	reg [7:0] programBufferMem_49;
	reg [7:0] programBufferMem_50;
	reg [7:0] programBufferMem_51;
	reg [7:0] programBufferMem_52;
	reg [7:0] programBufferMem_53;
	reg [7:0] programBufferMem_54;
	reg [7:0] programBufferMem_55;
	reg [7:0] programBufferMem_56;
	reg [7:0] programBufferMem_57;
	reg [7:0] programBufferMem_58;
	reg [7:0] programBufferMem_59;
	reg [7:0] programBufferMem_60;
	reg [7:0] programBufferMem_61;
	reg [7:0] programBufferMem_62;
	reg [7:0] programBufferMem_63;
	wire _resumeReqRegs_T = ~hartIsInResetSync_0;
	wire _resumeReqRegs_T_1 = resumeReqRegs & ~hartIsInResetSync_0;
	wire [1:0] _GEN_3655 = {1'd0, haltedBitRegs};
	wire [1:0] _haltedBitRegs_T = _GEN_3655 | 2'h1;
	wire [1:0] _GEN_3656 = {1'd0, _resumeReqRegs_T};
	wire [1:0] _haltedBitRegs_T_2 = _haltedBitRegs_T & _GEN_3656;
	wire [1:0] _haltedBitRegs_T_4 = _GEN_3655 & 2'h2;
	wire [1:0] _haltedBitRegs_T_6 = _haltedBitRegs_T_4 & _GEN_3656;
	wire _haltedBitRegs_T_8 = haltedBitRegs & _resumeReqRegs_T;
	wire out_backSel_66 = _out_backSel_T_1[66];
	wire out_woready_1_708 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_backSel_66) & (out_findex_1 == 10'h000);
	wire out_f_woready_808 = out_woready_1_708 & out_womask_941;
	wire [1:0] _GEN_61 = (out_f_woready_808 ? _haltedBitRegs_T_6 : {1'd0, _haltedBitRegs_T_8});
	wire out_backSel_64 = _out_backSel_T_1[64];
	wire out_woready_1_547 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_backSel_64) & (out_findex_1 == 10'h000);
	wire out_f_woready_647 = out_woready_1_547 & out_womask_941;
	wire [1:0] _GEN_62 = (out_f_woready_647 ? _haltedBitRegs_T_2 : _GEN_61);
	wire [1:0] _GEN_3659 = {1'd0, resumeReqRegs};
	wire [1:0] _resumeReqRegs_T_3 = _GEN_3659 & 2'h2;
	wire [1:0] _resumeReqRegs_T_5 = _resumeReqRegs_T_3 & _GEN_3656;
	wire [1:0] _GEN_63 = (out_f_woready_808 ? _resumeReqRegs_T_5 : {1'd0, _resumeReqRegs_T_1});
	wire _resumeReqRegs_T_8 = (resumeReqRegs | hamaskWrSel_0) & _resumeReqRegs_T;
	wire [1:0] _GEN_64 = (resumereq ? {1'd0, _resumeReqRegs_T_8} : _GEN_63);
	wire [1:0] _GEN_65 = (_T_1 ? 2'h0 : _GEN_62);
	wire [1:0] _GEN_66 = (_T_1 ? 2'h0 : _GEN_64);
	wire [31:0] out_prepend_2 = {programBufferMem_43, programBufferMem_42, programBufferMem_41, programBufferMem_40};
	wire [1:0] out_prepend_3 = {1'h0, ABSTRACTAUTOReg_autoexecdata[0]};
	wire [15:0] _out_T_108 = {14'd0, out_prepend_3};
	wire [31:0] out_prepend_4 = {ABSTRACTAUTOReg_autoexecprogbuf, _out_T_108};
	wire [31:0] out_prepend_7 = {programBufferMem_23, programBufferMem_22, programBufferMem_21, programBufferMem_20};
	wire [31:0] out_prepend_10 = {programBufferMem_59, programBufferMem_58, programBufferMem_57, programBufferMem_56};
	wire [31:0] out_prepend_13 = {programBufferMem_27, programBufferMem_26, programBufferMem_25, programBufferMem_24};
	wire [31:0] out_prepend_16 = {programBufferMem_7, programBufferMem_6, programBufferMem_5, programBufferMem_4};
	wire [31:0] out_prepend_19 = {programBufferMem_39, programBufferMem_38, programBufferMem_37, programBufferMem_36};
	wire [31:0] out_prepend_22 = {programBufferMem_3, programBufferMem_2, programBufferMem_1, programBufferMem_0};
	wire [31:0] out_prepend_25 = {programBufferMem_11, programBufferMem_10, programBufferMem_9, programBufferMem_8};
	wire [31:0] out_prepend_28 = {programBufferMem_55, programBufferMem_54, programBufferMem_53, programBufferMem_52};
	wire [16:0] out_prepend_41 = {resumeAcks, 1'h0, 1'h0, 1'h0, 1'h0, _T_10, _T_10, haltedBitRegs, haltedBitRegs, 8'ha2};
	wire [20:0] out_prepend_45 = {1'h0, haveResetBitRegs, haveResetBitRegs, resumeAcks, out_prepend_41};
	wire [21:0] _out_T_642 = {1'd0, out_prepend_45};
	wire [22:0] out_prepend_46 = {1'h0, _out_T_642};
	wire abstractCommandBusy = ctrlStateReg != 2'h0;
	wire [13:0] out_prepend_51 = {1'h0, abstractCommandBusy, 1'h0, ABSTRACTCSReg_cmderr, 8'h01};
	wire [23:0] _out_T_707 = {10'd0, out_prepend_51};
	wire [28:0] out_prepend_52 = {5'h10, _out_T_707};
	wire [31:0] out_prepend_55 = {programBufferMem_51, programBufferMem_50, programBufferMem_49, programBufferMem_48};
	wire [31:0] out_prepend_58 = {programBufferMem_31, programBufferMem_30, programBufferMem_29, programBufferMem_28};
	wire [31:0] out_prepend_61 = {programBufferMem_15, programBufferMem_14, programBufferMem_13, programBufferMem_12};
	wire [31:0] out_prepend_64 = {programBufferMem_47, programBufferMem_46, programBufferMem_45, programBufferMem_44};
	wire [31:0] out_prepend_67 = {programBufferMem_35, programBufferMem_34, programBufferMem_33, programBufferMem_32};
	wire [31:0] out_prepend_70 = {programBufferMem_19, programBufferMem_18, programBufferMem_17, programBufferMem_16};
	wire [31:0] out_prepend_73 = {abstractDataMem_3, abstractDataMem_2, abstractDataMem_1, abstractDataMem_0};
	wire [31:0] out_prepend_76 = {programBufferMem_63, programBufferMem_62, programBufferMem_61, programBufferMem_60};
	wire _GEN_266 = (5'h01 == out_iindex ? _out_T_2 : _out_T_20);
	wire _GEN_268 = (5'h03 == out_iindex ? _out_T_2 : (5'h02 == out_iindex) | _GEN_266);
	wire _GEN_269 = (5'h04 == out_iindex ? _out_T_44 : _GEN_268);
	wire _GEN_271 = (5'h06 == out_iindex ? _out_T_2 : (5'h05 == out_iindex) | _GEN_269);
	wire _GEN_272 = (5'h07 == out_iindex ? _out_T_2 : _GEN_271);
	wire _GEN_273 = (5'h08 == out_iindex ? _out_T_2 : _GEN_272);
	wire _GEN_281 = (5'h10 == out_iindex ? _out_T_44 : (5'h0f == out_iindex) | ((5'h0e == out_iindex) | ((5'h0d == out_iindex) | ((5'h0c == out_iindex) | ((5'h0b == out_iindex) | ((5'h0a == out_iindex) | ((5'h09 == out_iindex) | _GEN_273)))))));
	wire _GEN_282 = (5'h11 == out_iindex ? _out_T_44 : _GEN_281);
	wire _GEN_283 = (5'h12 == out_iindex ? _out_T_44 : _GEN_282);
	wire _GEN_284 = (5'h13 == out_iindex ? _out_T_44 : _GEN_283);
	wire _GEN_285 = (5'h14 == out_iindex ? _out_T_44 : _GEN_284);
	wire _GEN_286 = (5'h15 == out_iindex ? _out_T_44 : _GEN_285);
	wire _GEN_287 = (5'h16 == out_iindex ? _out_T_44 : _GEN_286);
	wire _GEN_288 = (5'h17 == out_iindex ? _out_T_44 : _GEN_287);
	wire _GEN_289 = (5'h18 == out_iindex ? _out_T_44 : _GEN_288);
	wire _GEN_290 = (5'h19 == out_iindex ? _out_T_44 : _GEN_289);
	wire _GEN_291 = (5'h1a == out_iindex ? _out_T_44 : _GEN_290);
	wire _GEN_292 = (5'h1b == out_iindex ? _out_T_44 : _GEN_291);
	wire _GEN_293 = (5'h1c == out_iindex ? _out_T_44 : _GEN_292);
	wire _GEN_294 = (5'h1d == out_iindex ? _out_T_44 : _GEN_293);
	wire _GEN_295 = (5'h1e == out_iindex ? _out_T_44 : _GEN_294);
	wire _GEN_296 = (5'h1f == out_iindex ? _out_T_44 : _GEN_295);
	wire [31:0] _out_out_bits_data_WIRE_1_1 = {9'd0, out_prepend_46};
	wire [31:0] _GEN_298 = (5'h01 == out_iindex ? _out_out_bits_data_WIRE_1_1 : haltedStatus_0);
	wire [31:0] _GEN_299 = (5'h02 == out_iindex ? 32'h00000000 : _GEN_298);
	wire [31:0] _GEN_300 = (5'h03 == out_iindex ? HALTSUM1RdData_haltsum1 : _GEN_299);
	wire [31:0] _GEN_301 = (5'h04 == out_iindex ? out_prepend_73 : _GEN_300);
	wire [31:0] _GEN_302 = (5'h05 == out_iindex ? 32'h00000000 : _GEN_301);
	wire [31:0] _out_out_bits_data_WIRE_1_6 = {3'd0, out_prepend_52};
	wire [31:0] _GEN_303 = (5'h06 == out_iindex ? _out_out_bits_data_WIRE_1_6 : _GEN_302);
	wire [31:0] _GEN_304 = (5'h07 == out_iindex ? _accessRegisterCommandReg_T : _GEN_303);
	wire [31:0] _GEN_305 = (5'h08 == out_iindex ? out_prepend_4 : _GEN_304);
	wire [31:0] _GEN_306 = (5'h09 == out_iindex ? 32'h00000000 : _GEN_305);
	wire [31:0] _GEN_307 = (5'h0a == out_iindex ? 32'h00000000 : _GEN_306);
	wire [31:0] _GEN_308 = (5'h0b == out_iindex ? 32'h00000000 : _GEN_307);
	wire [31:0] _GEN_309 = (5'h0c == out_iindex ? 32'h00000000 : _GEN_308);
	wire [31:0] _GEN_310 = (5'h0d == out_iindex ? 32'h00000000 : _GEN_309);
	wire [31:0] _GEN_311 = (5'h0e == out_iindex ? 32'h00000000 : _GEN_310);
	wire [31:0] _GEN_312 = (5'h0f == out_iindex ? 32'h00000000 : _GEN_311);
	wire [31:0] _GEN_313 = (5'h10 == out_iindex ? out_prepend_22 : _GEN_312);
	wire [31:0] _GEN_314 = (5'h11 == out_iindex ? out_prepend_16 : _GEN_313);
	wire [31:0] _GEN_315 = (5'h12 == out_iindex ? out_prepend_25 : _GEN_314);
	wire [31:0] _GEN_316 = (5'h13 == out_iindex ? out_prepend_61 : _GEN_315);
	wire [31:0] _GEN_317 = (5'h14 == out_iindex ? out_prepend_70 : _GEN_316);
	wire [31:0] _GEN_318 = (5'h15 == out_iindex ? out_prepend_7 : _GEN_317);
	wire [31:0] _GEN_319 = (5'h16 == out_iindex ? out_prepend_13 : _GEN_318);
	wire [31:0] _GEN_320 = (5'h17 == out_iindex ? out_prepend_58 : _GEN_319);
	wire [31:0] _GEN_321 = (5'h18 == out_iindex ? out_prepend_67 : _GEN_320);
	wire [31:0] _GEN_322 = (5'h19 == out_iindex ? out_prepend_19 : _GEN_321);
	wire [31:0] _GEN_323 = (5'h1a == out_iindex ? out_prepend_2 : _GEN_322);
	wire [31:0] _GEN_324 = (5'h1b == out_iindex ? out_prepend_64 : _GEN_323);
	wire [31:0] _GEN_325 = (5'h1c == out_iindex ? out_prepend_55 : _GEN_324);
	wire [31:0] _GEN_326 = (5'h1d == out_iindex ? out_prepend_28 : _GEN_325);
	wire [31:0] _GEN_327 = (5'h1e == out_iindex ? out_prepend_10 : _GEN_326);
	wire [31:0] _GEN_328 = (5'h1f == out_iindex ? out_prepend_76 : _GEN_327);
	reg goReg;
	wire [9:0] hartGoingId = auto_tl_in_a_bits_data[9:0];
	wire _T_341 = ~reset;
	wire _T_342 = ~(hartGoingId == 10'h000);
	wire out_backSel_65 = _out_backSel_T_1[65];
	wire out_woready_1_370 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_backSel_65) & (out_findex_1 == 10'h000);
	wire out_f_woready_470 = out_woready_1_370 & out_womask_941;
	wire _GEN_397 = (out_f_woready_470 ? 1'h0 : goReg);
	wire _GEN_3628 = (commandRegBadHaltResume ? 1'h0 : 1'h1);
	wire _GEN_3632 = (commandRegIsUnsupported ? 1'h0 : _GEN_3628);
	wire _GEN_3645 = (ctrlStateReg == 2'h1) & _GEN_3632;
	wire goAbstract = (ABSTRACTCSWrEnLegal ? 1'h0 : _GEN_3645);
	wire _GEN_398 = goAbstract | _GEN_397;
	wire accessRegisterCommandReg_postexec = _accessRegisterCommandReg_T[18];
	reg [31:0] abstractGeneratedMem_0;
	reg [31:0] abstractGeneratedMem_1;
	wire [15:0] _abstractGeneratedMem_0_inst_rd_T = accessRegisterCommandReg_regno & 16'h001f;
	wire [4:0] abstractGeneratedMem_0_inst_rd = _abstractGeneratedMem_0_inst_rd_T[4:0];
	wire [31:0] _abstractGeneratedMem_0_T = {17'h07000, accessRegisterCommandReg_size, abstractGeneratedMem_0_inst_rd, 7'h03};
	wire [31:0] _abstractGeneratedMem_0_T_1 = {7'h1c, abstractGeneratedMem_0_inst_rd, 5'h00, accessRegisterCommandReg_size, 5'h00, 7'h23};
	wire out_wimask_100 = &out_backMask_1[7:0];
	wire out_wimask_101 = &out_backMask_1[15:8];
	wire out_wimask_102 = &out_backMask_1[23:16];
	wire [23:0] out_prepend_78 = {6'h00, resumeReqRegs, goReg, 6'h00, resumeReqRegs, goReg, 6'h00, resumeReqRegs, goReg};
	wire out_wimask_103 = &out_backMask_1[31:24];
	wire [31:0] out_prepend_79 = {6'h00, resumeReqRegs, goReg, out_prepend_78};
	wire out_frontSel_217 = _out_backSel_T_1[217];
	wire out_wivalid_1_40 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_217) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_140 = out_wivalid_1_40 & out_wimask_100;
	wire out_f_wivalid_141 = out_wivalid_1_40 & out_wimask_101;
	wire out_f_wivalid_142 = out_wivalid_1_40 & out_wimask_102;
	wire out_f_wivalid_143 = out_wivalid_1_40 & out_wimask_103;
	wire out_frontSel_216 = _out_backSel_T_1[216];
	wire out_wivalid_1_176 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_216) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_276 = out_wivalid_1_176 & out_wimask_100;
	wire out_f_wivalid_277 = out_wivalid_1_176 & out_wimask_101;
	wire out_f_wivalid_278 = out_wivalid_1_176 & out_wimask_102;
	wire out_f_wivalid_279 = out_wivalid_1_176 & out_wimask_103;
	wire out_frontSel_211 = _out_backSel_T_1[211];
	wire out_wivalid_1_200 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_211) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_300 = out_wivalid_1_200 & out_wimask_100;
	wire out_f_wivalid_301 = out_wivalid_1_200 & out_wimask_101;
	wire out_f_wivalid_302 = out_wivalid_1_200 & out_wimask_102;
	wire out_f_wivalid_303 = out_wivalid_1_200 & out_wimask_103;
	wire out_frontSel_221 = _out_backSel_T_1[221];
	wire out_wivalid_1_232 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_221) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_332 = out_wivalid_1_232 & out_wimask_100;
	wire out_f_wivalid_333 = out_wivalid_1_232 & out_wimask_101;
	wire out_f_wivalid_334 = out_wivalid_1_232 & out_wimask_102;
	wire out_f_wivalid_335 = out_wivalid_1_232 & out_wimask_103;
	wire out_frontSel_220 = _out_backSel_T_1[220];
	wire out_wivalid_1_309 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_220) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_409 = out_wivalid_1_309 & out_wimask_100;
	wire out_f_wivalid_410 = out_wivalid_1_309 & out_wimask_101;
	wire out_f_wivalid_411 = out_wivalid_1_309 & out_wimask_102;
	wire out_f_wivalid_412 = out_wivalid_1_309 & out_wimask_103;
	wire out_frontSel_224 = _out_backSel_T_1[224];
	wire out_wivalid_1_403 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_224) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_503 = out_wivalid_1_403 & out_wimask_100;
	wire out_f_wivalid_504 = out_wivalid_1_403 & out_wimask_101;
	wire out_f_wivalid_505 = out_wivalid_1_403 & out_wimask_102;
	wire out_f_wivalid_506 = out_wivalid_1_403 & out_wimask_103;
	wire out_frontSel_212 = _out_backSel_T_1[212];
	wire out_wivalid_1_467 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_212) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_567 = out_wivalid_1_467 & out_wimask_100;
	wire out_f_wivalid_568 = out_wivalid_1_467 & out_wimask_101;
	wire out_f_wivalid_569 = out_wivalid_1_467 & out_wimask_102;
	wire out_f_wivalid_570 = out_wivalid_1_467 & out_wimask_103;
	wire out_frontSel_219 = _out_backSel_T_1[219];
	wire out_wivalid_1_624 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_219) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_724 = out_wivalid_1_624 & out_wimask_100;
	wire out_f_wivalid_725 = out_wivalid_1_624 & out_wimask_101;
	wire out_f_wivalid_726 = out_wivalid_1_624 & out_wimask_102;
	wire out_f_wivalid_727 = out_wivalid_1_624 & out_wimask_103;
	wire out_frontSel_208 = _out_backSel_T_1[208];
	wire out_wivalid_1_668 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_208) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_768 = out_wivalid_1_668 & out_wimask_100;
	wire out_f_wivalid_769 = out_wivalid_1_668 & out_wimask_101;
	wire out_f_wivalid_770 = out_wivalid_1_668 & out_wimask_102;
	wire out_f_wivalid_771 = out_wivalid_1_668 & out_wimask_103;
	wire out_frontSel_213 = _out_backSel_T_1[213];
	wire out_wivalid_1_696 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_213) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_796 = out_wivalid_1_696 & out_wimask_100;
	wire out_f_wivalid_797 = out_wivalid_1_696 & out_wimask_101;
	wire out_f_wivalid_798 = out_wivalid_1_696 & out_wimask_102;
	wire out_f_wivalid_799 = out_wivalid_1_696 & out_wimask_103;
	wire out_frontSel_223 = _out_backSel_T_1[223];
	wire out_wivalid_1_733 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_223) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_833 = out_wivalid_1_733 & out_wimask_100;
	wire out_f_wivalid_834 = out_wivalid_1_733 & out_wimask_101;
	wire out_f_wivalid_835 = out_wivalid_1_733 & out_wimask_102;
	wire out_f_wivalid_836 = out_wivalid_1_733 & out_wimask_103;
	wire out_frontSel_209 = _out_backSel_T_1[209];
	wire out_wivalid_1_785 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_209) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_885 = out_wivalid_1_785 & out_wimask_100;
	wire out_f_wivalid_886 = out_wivalid_1_785 & out_wimask_101;
	wire out_f_wivalid_887 = out_wivalid_1_785 & out_wimask_102;
	wire out_f_wivalid_888 = out_wivalid_1_785 & out_wimask_103;
	wire out_frontSel_218 = _out_backSel_T_1[218];
	wire out_wivalid_1_918 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_218) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_1018 = out_wivalid_1_918 & out_wimask_100;
	wire out_f_wivalid_1019 = out_wivalid_1_918 & out_wimask_101;
	wire out_f_wivalid_1020 = out_wivalid_1_918 & out_wimask_102;
	wire out_f_wivalid_1021 = out_wivalid_1_918 & out_wimask_103;
	wire out_frontSel_214 = _out_backSel_T_1[214];
	wire out_wivalid_1_991 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_214) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_1091 = out_wivalid_1_991 & out_wimask_100;
	wire out_f_wivalid_1092 = out_wivalid_1_991 & out_wimask_101;
	wire out_f_wivalid_1093 = out_wivalid_1_991 & out_wimask_102;
	wire out_f_wivalid_1094 = out_wivalid_1_991 & out_wimask_103;
	wire out_frontSel_210 = _out_backSel_T_1[210];
	wire out_wivalid_1_1043 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_210) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_1143 = out_wivalid_1_1043 & out_wimask_100;
	wire out_f_wivalid_1144 = out_wivalid_1_1043 & out_wimask_101;
	wire out_f_wivalid_1145 = out_wivalid_1_1043 & out_wimask_102;
	wire out_f_wivalid_1146 = out_wivalid_1_1043 & out_wimask_103;
	wire out_frontSel_215 = _out_backSel_T_1[215];
	wire out_wivalid_1_1159 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_215) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_1259 = out_wivalid_1_1159 & out_wimask_100;
	wire out_f_wivalid_1260 = out_wivalid_1_1159 & out_wimask_101;
	wire out_f_wivalid_1261 = out_wivalid_1_1159 & out_wimask_102;
	wire out_f_wivalid_1262 = out_wivalid_1_1159 & out_wimask_103;
	wire out_frontSel_222 = _out_backSel_T_1[222];
	wire out_wivalid_1_1167 = (((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_1_bits_read) & out_frontSel_222) & (out_findex_1 == 10'h000);
	wire out_f_wivalid_1267 = out_wivalid_1_1167 & out_wimask_100;
	wire out_f_wivalid_1268 = out_wivalid_1_1167 & out_wimask_101;
	wire out_f_wivalid_1269 = out_wivalid_1_1167 & out_wimask_102;
	wire out_f_wivalid_1270 = out_wivalid_1_1167 & out_wimask_103;
	wire _GEN_2523 = (9'h001 == out_iindex_1 ? _out_T_1642 : _out_T_1642);
	wire _GEN_2524 = (9'h002 == out_iindex_1 ? _out_T_1642 : _GEN_2523);
	wire _GEN_2525 = (9'h003 == out_iindex_1 ? _out_T_1642 : _GEN_2524);
	wire _GEN_2526 = (9'h004 == out_iindex_1 ? _out_T_1642 : _GEN_2525);
	wire _GEN_2527 = (9'h005 == out_iindex_1 ? _out_T_1642 : _GEN_2526);
	wire _GEN_2528 = (9'h006 == out_iindex_1 ? _out_T_1642 : _GEN_2527);
	wire _GEN_2529 = (9'h007 == out_iindex_1 ? _out_T_1642 : _GEN_2528);
	wire _GEN_2530 = (9'h008 == out_iindex_1 ? _out_T_1642 : _GEN_2529);
	wire _GEN_2531 = (9'h009 == out_iindex_1 ? _out_T_1642 : _GEN_2530);
	wire _GEN_2532 = (9'h00a == out_iindex_1 ? _out_T_1642 : _GEN_2531);
	wire _GEN_2533 = (9'h00b == out_iindex_1 ? _out_T_1642 : _GEN_2532);
	wire _GEN_2534 = (9'h00c == out_iindex_1 ? _out_T_1642 : _GEN_2533);
	wire _GEN_2535 = (9'h00d == out_iindex_1 ? _out_T_1642 : _GEN_2534);
	wire _GEN_2536 = (9'h00e == out_iindex_1 ? _out_T_1642 : _GEN_2535);
	wire _GEN_2537 = (9'h00f == out_iindex_1 ? _out_T_1642 : _GEN_2536);
	wire _GEN_2538 = (9'h010 == out_iindex_1 ? _out_T_1642 : _GEN_2537);
	wire _GEN_2539 = (9'h011 == out_iindex_1 ? _out_T_1642 : _GEN_2538);
	wire _GEN_2540 = (9'h012 == out_iindex_1 ? _out_T_1642 : _GEN_2539);
	wire _GEN_2541 = (9'h013 == out_iindex_1 ? _out_T_1642 : _GEN_2540);
	wire _GEN_2542 = (9'h014 == out_iindex_1 ? _out_T_1642 : _GEN_2541);
	wire _GEN_2557 = (9'h023 == out_iindex_1) | ((9'h022 == out_iindex_1) | ((9'h021 == out_iindex_1) | ((9'h020 == out_iindex_1) | ((9'h01f == out_iindex_1) | ((9'h01e == out_iindex_1) | ((9'h01d == out_iindex_1) | ((9'h01c == out_iindex_1) | ((9'h01b == out_iindex_1) | ((9'h01a == out_iindex_1) | ((9'h019 == out_iindex_1) | ((9'h018 == out_iindex_1) | ((9'h017 == out_iindex_1) | ((9'h016 == out_iindex_1) | ((9'h015 == out_iindex_1) | _GEN_2542))))))))))))));
	wire _GEN_2572 = (9'h032 == out_iindex_1) | ((9'h031 == out_iindex_1) | ((9'h030 == out_iindex_1) | ((9'h02f == out_iindex_1) | ((9'h02e == out_iindex_1) | ((9'h02d == out_iindex_1) | ((9'h02c == out_iindex_1) | ((9'h02b == out_iindex_1) | ((9'h02a == out_iindex_1) | ((9'h029 == out_iindex_1) | ((9'h028 == out_iindex_1) | ((9'h027 == out_iindex_1) | ((9'h026 == out_iindex_1) | ((9'h025 == out_iindex_1) | ((9'h024 == out_iindex_1) | _GEN_2557))))))))))))));
	wire _GEN_2586 = (9'h040 == out_iindex_1 ? _out_T_1122 : (9'h03f == out_iindex_1) | ((9'h03e == out_iindex_1) | ((9'h03d == out_iindex_1) | ((9'h03c == out_iindex_1) | ((9'h03b == out_iindex_1) | ((9'h03a == out_iindex_1) | ((9'h039 == out_iindex_1) | ((9'h038 == out_iindex_1) | ((9'h037 == out_iindex_1) | ((9'h036 == out_iindex_1) | ((9'h035 == out_iindex_1) | ((9'h034 == out_iindex_1) | ((9'h033 == out_iindex_1) | _GEN_2572)))))))))))));
	wire _GEN_2587 = (9'h041 == out_iindex_1 ? _out_T_1122 : _GEN_2586);
	wire _GEN_2588 = (9'h042 == out_iindex_1 ? _out_T_1122 : _GEN_2587);
	wire _GEN_2589 = (9'h043 == out_iindex_1 ? _out_T_1122 : _GEN_2588);
	wire _GEN_2604 = (9'h052 == out_iindex_1) | ((9'h051 == out_iindex_1) | ((9'h050 == out_iindex_1) | ((9'h04f == out_iindex_1) | ((9'h04e == out_iindex_1) | ((9'h04d == out_iindex_1) | ((9'h04c == out_iindex_1) | ((9'h04b == out_iindex_1) | ((9'h04a == out_iindex_1) | ((9'h049 == out_iindex_1) | ((9'h048 == out_iindex_1) | ((9'h047 == out_iindex_1) | ((9'h046 == out_iindex_1) | ((9'h045 == out_iindex_1) | ((9'h044 == out_iindex_1) | _GEN_2589))))))))))))));
	wire _GEN_2619 = (9'h061 == out_iindex_1) | ((9'h060 == out_iindex_1) | ((9'h05f == out_iindex_1) | ((9'h05e == out_iindex_1) | ((9'h05d == out_iindex_1) | ((9'h05c == out_iindex_1) | ((9'h05b == out_iindex_1) | ((9'h05a == out_iindex_1) | ((9'h059 == out_iindex_1) | ((9'h058 == out_iindex_1) | ((9'h057 == out_iindex_1) | ((9'h056 == out_iindex_1) | ((9'h055 == out_iindex_1) | ((9'h054 == out_iindex_1) | ((9'h053 == out_iindex_1) | _GEN_2604))))))))))))));
	wire _GEN_2634 = (9'h070 == out_iindex_1) | ((9'h06f == out_iindex_1) | ((9'h06e == out_iindex_1) | ((9'h06d == out_iindex_1) | ((9'h06c == out_iindex_1) | ((9'h06b == out_iindex_1) | ((9'h06a == out_iindex_1) | ((9'h069 == out_iindex_1) | ((9'h068 == out_iindex_1) | ((9'h067 == out_iindex_1) | ((9'h066 == out_iindex_1) | ((9'h065 == out_iindex_1) | ((9'h064 == out_iindex_1) | ((9'h063 == out_iindex_1) | ((9'h062 == out_iindex_1) | _GEN_2619))))))))))))));
	wire _GEN_2649 = (9'h07f == out_iindex_1) | ((9'h07e == out_iindex_1) | ((9'h07d == out_iindex_1) | ((9'h07c == out_iindex_1) | ((9'h07b == out_iindex_1) | ((9'h07a == out_iindex_1) | ((9'h079 == out_iindex_1) | ((9'h078 == out_iindex_1) | ((9'h077 == out_iindex_1) | ((9'h076 == out_iindex_1) | ((9'h075 == out_iindex_1) | ((9'h074 == out_iindex_1) | ((9'h073 == out_iindex_1) | ((9'h072 == out_iindex_1) | ((9'h071 == out_iindex_1) | _GEN_2634))))))))))))));
	wire _GEN_2664 = (9'h08e == out_iindex_1) | ((9'h08d == out_iindex_1) | ((9'h08c == out_iindex_1) | ((9'h08b == out_iindex_1) | ((9'h08a == out_iindex_1) | ((9'h089 == out_iindex_1) | ((9'h088 == out_iindex_1) | ((9'h087 == out_iindex_1) | ((9'h086 == out_iindex_1) | ((9'h085 == out_iindex_1) | ((9'h084 == out_iindex_1) | ((9'h083 == out_iindex_1) | ((9'h082 == out_iindex_1) | ((9'h081 == out_iindex_1) | ((9'h080 == out_iindex_1) | _GEN_2649))))))))))))));
	wire _GEN_2679 = (9'h09d == out_iindex_1) | ((9'h09c == out_iindex_1) | ((9'h09b == out_iindex_1) | ((9'h09a == out_iindex_1) | ((9'h099 == out_iindex_1) | ((9'h098 == out_iindex_1) | ((9'h097 == out_iindex_1) | ((9'h096 == out_iindex_1) | ((9'h095 == out_iindex_1) | ((9'h094 == out_iindex_1) | ((9'h093 == out_iindex_1) | ((9'h092 == out_iindex_1) | ((9'h091 == out_iindex_1) | ((9'h090 == out_iindex_1) | ((9'h08f == out_iindex_1) | _GEN_2664))))))))))))));
	wire _GEN_2694 = (9'h0ac == out_iindex_1) | ((9'h0ab == out_iindex_1) | ((9'h0aa == out_iindex_1) | ((9'h0a9 == out_iindex_1) | ((9'h0a8 == out_iindex_1) | ((9'h0a7 == out_iindex_1) | ((9'h0a6 == out_iindex_1) | ((9'h0a5 == out_iindex_1) | ((9'h0a4 == out_iindex_1) | ((9'h0a3 == out_iindex_1) | ((9'h0a2 == out_iindex_1) | ((9'h0a1 == out_iindex_1) | ((9'h0a0 == out_iindex_1) | ((9'h09f == out_iindex_1) | ((9'h09e == out_iindex_1) | _GEN_2679))))))))))))));
	wire _GEN_2709 = (9'h0bb == out_iindex_1) | ((9'h0ba == out_iindex_1) | ((9'h0b9 == out_iindex_1) | ((9'h0b8 == out_iindex_1) | ((9'h0b7 == out_iindex_1) | ((9'h0b6 == out_iindex_1) | ((9'h0b5 == out_iindex_1) | ((9'h0b4 == out_iindex_1) | ((9'h0b3 == out_iindex_1) | ((9'h0b2 == out_iindex_1) | ((9'h0b1 == out_iindex_1) | ((9'h0b0 == out_iindex_1) | ((9'h0af == out_iindex_1) | ((9'h0ae == out_iindex_1) | ((9'h0ad == out_iindex_1) | _GEN_2694))))))))))))));
	wire _GEN_2714 = (9'h0c0 == out_iindex_1 ? _out_T_1122 : (9'h0bf == out_iindex_1) | ((9'h0be == out_iindex_1) | ((9'h0bd == out_iindex_1) | ((9'h0bc == out_iindex_1) | _GEN_2709))));
	wire _GEN_2728 = (9'h0ce == out_iindex_1 ? _out_T_1122 : (9'h0cd == out_iindex_1) | ((9'h0cc == out_iindex_1) | ((9'h0cb == out_iindex_1) | ((9'h0ca == out_iindex_1) | ((9'h0c9 == out_iindex_1) | ((9'h0c8 == out_iindex_1) | ((9'h0c7 == out_iindex_1) | ((9'h0c6 == out_iindex_1) | ((9'h0c5 == out_iindex_1) | ((9'h0c4 == out_iindex_1) | ((9'h0c3 == out_iindex_1) | ((9'h0c2 == out_iindex_1) | ((9'h0c1 == out_iindex_1) | _GEN_2714)))))))))))));
	wire _GEN_2729 = (9'h0cf == out_iindex_1 ? _out_T_1122 : _GEN_2728);
	wire _GEN_2730 = (9'h0d0 == out_iindex_1 ? _out_T_1122 : _GEN_2729);
	wire _GEN_2731 = (9'h0d1 == out_iindex_1 ? _out_T_1122 : _GEN_2730);
	wire _GEN_2732 = (9'h0d2 == out_iindex_1 ? _out_T_1122 : _GEN_2731);
	wire _GEN_2733 = (9'h0d3 == out_iindex_1 ? _out_T_1122 : _GEN_2732);
	wire _GEN_2734 = (9'h0d4 == out_iindex_1 ? _out_T_1122 : _GEN_2733);
	wire _GEN_2735 = (9'h0d5 == out_iindex_1 ? _out_T_1122 : _GEN_2734);
	wire _GEN_2736 = (9'h0d6 == out_iindex_1 ? _out_T_1122 : _GEN_2735);
	wire _GEN_2737 = (9'h0d7 == out_iindex_1 ? _out_T_1122 : _GEN_2736);
	wire _GEN_2738 = (9'h0d8 == out_iindex_1 ? _out_T_1122 : _GEN_2737);
	wire _GEN_2739 = (9'h0d9 == out_iindex_1 ? _out_T_1122 : _GEN_2738);
	wire _GEN_2740 = (9'h0da == out_iindex_1 ? _out_T_1122 : _GEN_2739);
	wire _GEN_2741 = (9'h0db == out_iindex_1 ? _out_T_1122 : _GEN_2740);
	wire _GEN_2742 = (9'h0dc == out_iindex_1 ? _out_T_1122 : _GEN_2741);
	wire _GEN_2743 = (9'h0dd == out_iindex_1 ? _out_T_1122 : _GEN_2742);
	wire _GEN_2744 = (9'h0de == out_iindex_1 ? _out_T_1122 : _GEN_2743);
	wire _GEN_2745 = (9'h0df == out_iindex_1 ? _out_T_1122 : _GEN_2744);
	wire _GEN_2746 = (9'h0e0 == out_iindex_1 ? _out_T_1122 : _GEN_2745);
	wire _GEN_2761 = (9'h0ef == out_iindex_1) | ((9'h0ee == out_iindex_1) | ((9'h0ed == out_iindex_1) | ((9'h0ec == out_iindex_1) | ((9'h0eb == out_iindex_1) | ((9'h0ea == out_iindex_1) | ((9'h0e9 == out_iindex_1) | ((9'h0e8 == out_iindex_1) | ((9'h0e7 == out_iindex_1) | ((9'h0e6 == out_iindex_1) | ((9'h0e5 == out_iindex_1) | ((9'h0e4 == out_iindex_1) | ((9'h0e3 == out_iindex_1) | ((9'h0e2 == out_iindex_1) | ((9'h0e1 == out_iindex_1) | _GEN_2746))))))))))))));
	wire _GEN_2776 = (9'h0fe == out_iindex_1) | ((9'h0fd == out_iindex_1) | ((9'h0fc == out_iindex_1) | ((9'h0fb == out_iindex_1) | ((9'h0fa == out_iindex_1) | ((9'h0f9 == out_iindex_1) | ((9'h0f8 == out_iindex_1) | ((9'h0f7 == out_iindex_1) | ((9'h0f6 == out_iindex_1) | ((9'h0f5 == out_iindex_1) | ((9'h0f4 == out_iindex_1) | ((9'h0f3 == out_iindex_1) | ((9'h0f2 == out_iindex_1) | ((9'h0f1 == out_iindex_1) | ((9'h0f0 == out_iindex_1) | _GEN_2761))))))))))))));
	wire _GEN_2778 = (9'h100 == out_iindex_1 ? _out_T_1122 : (9'h0ff == out_iindex_1) | _GEN_2776);
	wire _GEN_2779 = (9'h101 == out_iindex_1 ? _out_T_1122 : _GEN_2778);
	wire _GEN_2780 = (9'h102 == out_iindex_1 ? _out_T_1122 : _GEN_2779);
	wire _GEN_2781 = (9'h103 == out_iindex_1 ? _out_T_1122 : _GEN_2780);
	wire _GEN_2782 = (9'h104 == out_iindex_1 ? _out_T_1122 : _GEN_2781);
	wire _GEN_2783 = (9'h105 == out_iindex_1 ? _out_T_1122 : _GEN_2782);
	wire _GEN_2784 = (9'h106 == out_iindex_1 ? _out_T_1122 : _GEN_2783);
	wire _GEN_2785 = (9'h107 == out_iindex_1 ? _out_T_1122 : _GEN_2784);
	wire _GEN_2786 = (9'h108 == out_iindex_1 ? _out_T_1122 : _GEN_2785);
	wire _GEN_2787 = (9'h109 == out_iindex_1 ? _out_T_1122 : _GEN_2786);
	wire _GEN_2788 = (9'h10a == out_iindex_1 ? _out_T_1122 : _GEN_2787);
	wire _GEN_2789 = (9'h10b == out_iindex_1 ? _out_T_1122 : _GEN_2788);
	wire _GEN_2790 = (9'h10c == out_iindex_1 ? _out_T_1122 : _GEN_2789);
	wire _GEN_2791 = (9'h10d == out_iindex_1 ? _out_T_1122 : _GEN_2790);
	wire _GEN_2792 = (9'h10e == out_iindex_1 ? _out_T_1122 : _GEN_2791);
	wire _GEN_2793 = (9'h10f == out_iindex_1 ? _out_T_1122 : _GEN_2792);
	wire _GEN_2794 = (9'h110 == out_iindex_1 ? _out_T_1122 : _GEN_2793);
	wire _GEN_2795 = (9'h111 == out_iindex_1 ? _out_T_1122 : _GEN_2794);
	wire _GEN_2796 = (9'h112 == out_iindex_1 ? _out_T_1122 : _GEN_2795);
	wire _GEN_2797 = (9'h113 == out_iindex_1 ? _out_T_1122 : _GEN_2796);
	wire _GEN_2798 = (9'h114 == out_iindex_1 ? _out_T_1122 : _GEN_2797);
	wire _GEN_2799 = (9'h115 == out_iindex_1 ? _out_T_1122 : _GEN_2798);
	wire _GEN_2800 = (9'h116 == out_iindex_1 ? _out_T_1122 : _GEN_2799);
	wire _GEN_2801 = (9'h117 == out_iindex_1 ? _out_T_1122 : _GEN_2800);
	wire _GEN_2802 = (9'h118 == out_iindex_1 ? _out_T_1122 : _GEN_2801);
	wire _GEN_2803 = (9'h119 == out_iindex_1 ? _out_T_1122 : _GEN_2802);
	wire _GEN_2804 = (9'h11a == out_iindex_1 ? _out_T_1122 : _GEN_2803);
	wire _GEN_2805 = (9'h11b == out_iindex_1 ? _out_T_1122 : _GEN_2804);
	wire _GEN_2806 = (9'h11c == out_iindex_1 ? _out_T_1122 : _GEN_2805);
	wire _GEN_2807 = (9'h11d == out_iindex_1 ? _out_T_1122 : _GEN_2806);
	wire _GEN_2808 = (9'h11e == out_iindex_1 ? _out_T_1122 : _GEN_2807);
	wire _GEN_2809 = (9'h11f == out_iindex_1 ? _out_T_1122 : _GEN_2808);
	wire _GEN_2810 = (9'h120 == out_iindex_1 ? _out_T_1122 : _GEN_2809);
	wire _GEN_2811 = (9'h121 == out_iindex_1 ? _out_T_1122 : _GEN_2810);
	wire _GEN_2812 = (9'h122 == out_iindex_1 ? _out_T_1122 : _GEN_2811);
	wire _GEN_2813 = (9'h123 == out_iindex_1 ? _out_T_1122 : _GEN_2812);
	wire _GEN_2814 = (9'h124 == out_iindex_1 ? _out_T_1122 : _GEN_2813);
	wire _GEN_2815 = (9'h125 == out_iindex_1 ? _out_T_1122 : _GEN_2814);
	wire _GEN_2816 = (9'h126 == out_iindex_1 ? _out_T_1122 : _GEN_2815);
	wire _GEN_2817 = (9'h127 == out_iindex_1 ? _out_T_1122 : _GEN_2816);
	wire _GEN_2818 = (9'h128 == out_iindex_1 ? _out_T_1122 : _GEN_2817);
	wire _GEN_2819 = (9'h129 == out_iindex_1 ? _out_T_1122 : _GEN_2818);
	wire _GEN_2820 = (9'h12a == out_iindex_1 ? _out_T_1122 : _GEN_2819);
	wire _GEN_2821 = (9'h12b == out_iindex_1 ? _out_T_1122 : _GEN_2820);
	wire _GEN_2822 = (9'h12c == out_iindex_1 ? _out_T_1122 : _GEN_2821);
	wire _GEN_2823 = (9'h12d == out_iindex_1 ? _out_T_1122 : _GEN_2822);
	wire _GEN_2824 = (9'h12e == out_iindex_1 ? _out_T_1122 : _GEN_2823);
	wire _GEN_2825 = (9'h12f == out_iindex_1 ? _out_T_1122 : _GEN_2824);
	wire _GEN_2826 = (9'h130 == out_iindex_1 ? _out_T_1122 : _GEN_2825);
	wire _GEN_2827 = (9'h131 == out_iindex_1 ? _out_T_1122 : _GEN_2826);
	wire _GEN_2828 = (9'h132 == out_iindex_1 ? _out_T_1122 : _GEN_2827);
	wire _GEN_2829 = (9'h133 == out_iindex_1 ? _out_T_1122 : _GEN_2828);
	wire _GEN_2830 = (9'h134 == out_iindex_1 ? _out_T_1122 : _GEN_2829);
	wire _GEN_2831 = (9'h135 == out_iindex_1 ? _out_T_1122 : _GEN_2830);
	wire _GEN_2832 = (9'h136 == out_iindex_1 ? _out_T_1122 : _GEN_2831);
	wire _GEN_2833 = (9'h137 == out_iindex_1 ? _out_T_1122 : _GEN_2832);
	wire _GEN_2834 = (9'h138 == out_iindex_1 ? _out_T_1122 : _GEN_2833);
	wire _GEN_2835 = (9'h139 == out_iindex_1 ? _out_T_1122 : _GEN_2834);
	wire _GEN_2836 = (9'h13a == out_iindex_1 ? _out_T_1122 : _GEN_2835);
	wire _GEN_2837 = (9'h13b == out_iindex_1 ? _out_T_1122 : _GEN_2836);
	wire _GEN_2838 = (9'h13c == out_iindex_1 ? _out_T_1122 : _GEN_2837);
	wire _GEN_2839 = (9'h13d == out_iindex_1 ? _out_T_1122 : _GEN_2838);
	wire _GEN_2840 = (9'h13e == out_iindex_1 ? _out_T_1122 : _GEN_2839);
	wire _GEN_2841 = (9'h13f == out_iindex_1 ? _out_T_1122 : _GEN_2840);
	wire _GEN_2842 = (9'h140 == out_iindex_1 ? _out_T_1122 : _GEN_2841);
	wire _GEN_2843 = (9'h141 == out_iindex_1 ? _out_T_1122 : _GEN_2842);
	wire _GEN_2844 = (9'h142 == out_iindex_1 ? _out_T_1122 : _GEN_2843);
	wire _GEN_2845 = (9'h143 == out_iindex_1 ? _out_T_1122 : _GEN_2844);
	wire _GEN_2846 = (9'h144 == out_iindex_1 ? _out_T_1122 : _GEN_2845);
	wire _GEN_2847 = (9'h145 == out_iindex_1 ? _out_T_1122 : _GEN_2846);
	wire _GEN_2848 = (9'h146 == out_iindex_1 ? _out_T_1122 : _GEN_2847);
	wire _GEN_2849 = (9'h147 == out_iindex_1 ? _out_T_1122 : _GEN_2848);
	wire _GEN_2850 = (9'h148 == out_iindex_1 ? _out_T_1122 : _GEN_2849);
	wire _GEN_2851 = (9'h149 == out_iindex_1 ? _out_T_1122 : _GEN_2850);
	wire _GEN_2852 = (9'h14a == out_iindex_1 ? _out_T_1122 : _GEN_2851);
	wire _GEN_2853 = (9'h14b == out_iindex_1 ? _out_T_1122 : _GEN_2852);
	wire _GEN_2854 = (9'h14c == out_iindex_1 ? _out_T_1122 : _GEN_2853);
	wire _GEN_2855 = (9'h14d == out_iindex_1 ? _out_T_1122 : _GEN_2854);
	wire _GEN_2856 = (9'h14e == out_iindex_1 ? _out_T_1122 : _GEN_2855);
	wire _GEN_2857 = (9'h14f == out_iindex_1 ? _out_T_1122 : _GEN_2856);
	wire _GEN_2858 = (9'h150 == out_iindex_1 ? _out_T_1122 : _GEN_2857);
	wire _GEN_2859 = (9'h151 == out_iindex_1 ? _out_T_1122 : _GEN_2858);
	wire _GEN_2860 = (9'h152 == out_iindex_1 ? _out_T_1122 : _GEN_2859);
	wire _GEN_2861 = (9'h153 == out_iindex_1 ? _out_T_1122 : _GEN_2860);
	wire _GEN_2862 = (9'h154 == out_iindex_1 ? _out_T_1122 : _GEN_2861);
	wire _GEN_2863 = (9'h155 == out_iindex_1 ? _out_T_1122 : _GEN_2862);
	wire _GEN_2864 = (9'h156 == out_iindex_1 ? _out_T_1122 : _GEN_2863);
	wire _GEN_2865 = (9'h157 == out_iindex_1 ? _out_T_1122 : _GEN_2864);
	wire _GEN_2866 = (9'h158 == out_iindex_1 ? _out_T_1122 : _GEN_2865);
	wire _GEN_2867 = (9'h159 == out_iindex_1 ? _out_T_1122 : _GEN_2866);
	wire _GEN_2868 = (9'h15a == out_iindex_1 ? _out_T_1122 : _GEN_2867);
	wire _GEN_2869 = (9'h15b == out_iindex_1 ? _out_T_1122 : _GEN_2868);
	wire _GEN_2870 = (9'h15c == out_iindex_1 ? _out_T_1122 : _GEN_2869);
	wire _GEN_2871 = (9'h15d == out_iindex_1 ? _out_T_1122 : _GEN_2870);
	wire _GEN_2872 = (9'h15e == out_iindex_1 ? _out_T_1122 : _GEN_2871);
	wire _GEN_2873 = (9'h15f == out_iindex_1 ? _out_T_1122 : _GEN_2872);
	wire _GEN_2874 = (9'h160 == out_iindex_1 ? _out_T_1122 : _GEN_2873);
	wire _GEN_2875 = (9'h161 == out_iindex_1 ? _out_T_1122 : _GEN_2874);
	wire _GEN_2876 = (9'h162 == out_iindex_1 ? _out_T_1122 : _GEN_2875);
	wire _GEN_2877 = (9'h163 == out_iindex_1 ? _out_T_1122 : _GEN_2876);
	wire _GEN_2878 = (9'h164 == out_iindex_1 ? _out_T_1122 : _GEN_2877);
	wire _GEN_2879 = (9'h165 == out_iindex_1 ? _out_T_1122 : _GEN_2878);
	wire _GEN_2880 = (9'h166 == out_iindex_1 ? _out_T_1122 : _GEN_2879);
	wire _GEN_2881 = (9'h167 == out_iindex_1 ? _out_T_1122 : _GEN_2880);
	wire _GEN_2882 = (9'h168 == out_iindex_1 ? _out_T_1122 : _GEN_2881);
	wire _GEN_2883 = (9'h169 == out_iindex_1 ? _out_T_1122 : _GEN_2882);
	wire _GEN_2884 = (9'h16a == out_iindex_1 ? _out_T_1122 : _GEN_2883);
	wire _GEN_2885 = (9'h16b == out_iindex_1 ? _out_T_1122 : _GEN_2884);
	wire _GEN_2886 = (9'h16c == out_iindex_1 ? _out_T_1122 : _GEN_2885);
	wire _GEN_2887 = (9'h16d == out_iindex_1 ? _out_T_1122 : _GEN_2886);
	wire _GEN_2888 = (9'h16e == out_iindex_1 ? _out_T_1122 : _GEN_2887);
	wire _GEN_2889 = (9'h16f == out_iindex_1 ? _out_T_1122 : _GEN_2888);
	wire _GEN_2890 = (9'h170 == out_iindex_1 ? _out_T_1122 : _GEN_2889);
	wire _GEN_2891 = (9'h171 == out_iindex_1 ? _out_T_1122 : _GEN_2890);
	wire _GEN_2892 = (9'h172 == out_iindex_1 ? _out_T_1122 : _GEN_2891);
	wire _GEN_2893 = (9'h173 == out_iindex_1 ? _out_T_1122 : _GEN_2892);
	wire _GEN_2894 = (9'h174 == out_iindex_1 ? _out_T_1122 : _GEN_2893);
	wire _GEN_2895 = (9'h175 == out_iindex_1 ? _out_T_1122 : _GEN_2894);
	wire _GEN_2896 = (9'h176 == out_iindex_1 ? _out_T_1122 : _GEN_2895);
	wire _GEN_2897 = (9'h177 == out_iindex_1 ? _out_T_1122 : _GEN_2896);
	wire _GEN_2898 = (9'h178 == out_iindex_1 ? _out_T_1122 : _GEN_2897);
	wire _GEN_2899 = (9'h179 == out_iindex_1 ? _out_T_1122 : _GEN_2898);
	wire _GEN_2900 = (9'h17a == out_iindex_1 ? _out_T_1122 : _GEN_2899);
	wire _GEN_2901 = (9'h17b == out_iindex_1 ? _out_T_1122 : _GEN_2900);
	wire _GEN_2902 = (9'h17c == out_iindex_1 ? _out_T_1122 : _GEN_2901);
	wire _GEN_2903 = (9'h17d == out_iindex_1 ? _out_T_1122 : _GEN_2902);
	wire _GEN_2904 = (9'h17e == out_iindex_1 ? _out_T_1122 : _GEN_2903);
	wire _GEN_2905 = (9'h17f == out_iindex_1 ? _out_T_1122 : _GEN_2904);
	wire _GEN_2906 = (9'h180 == out_iindex_1 ? _out_T_1122 : _GEN_2905);
	wire _GEN_2907 = (9'h181 == out_iindex_1 ? _out_T_1122 : _GEN_2906);
	wire _GEN_2908 = (9'h182 == out_iindex_1 ? _out_T_1122 : _GEN_2907);
	wire _GEN_2909 = (9'h183 == out_iindex_1 ? _out_T_1122 : _GEN_2908);
	wire _GEN_2910 = (9'h184 == out_iindex_1 ? _out_T_1122 : _GEN_2909);
	wire _GEN_2911 = (9'h185 == out_iindex_1 ? _out_T_1122 : _GEN_2910);
	wire _GEN_2912 = (9'h186 == out_iindex_1 ? _out_T_1122 : _GEN_2911);
	wire _GEN_2913 = (9'h187 == out_iindex_1 ? _out_T_1122 : _GEN_2912);
	wire _GEN_2914 = (9'h188 == out_iindex_1 ? _out_T_1122 : _GEN_2913);
	wire _GEN_2915 = (9'h189 == out_iindex_1 ? _out_T_1122 : _GEN_2914);
	wire _GEN_2916 = (9'h18a == out_iindex_1 ? _out_T_1122 : _GEN_2915);
	wire _GEN_2917 = (9'h18b == out_iindex_1 ? _out_T_1122 : _GEN_2916);
	wire _GEN_2918 = (9'h18c == out_iindex_1 ? _out_T_1122 : _GEN_2917);
	wire _GEN_2919 = (9'h18d == out_iindex_1 ? _out_T_1122 : _GEN_2918);
	wire _GEN_2920 = (9'h18e == out_iindex_1 ? _out_T_1122 : _GEN_2919);
	wire _GEN_2921 = (9'h18f == out_iindex_1 ? _out_T_1122 : _GEN_2920);
	wire _GEN_2922 = (9'h190 == out_iindex_1 ? _out_T_1122 : _GEN_2921);
	wire _GEN_2923 = (9'h191 == out_iindex_1 ? _out_T_1122 : _GEN_2922);
	wire _GEN_2924 = (9'h192 == out_iindex_1 ? _out_T_1122 : _GEN_2923);
	wire _GEN_2925 = (9'h193 == out_iindex_1 ? _out_T_1122 : _GEN_2924);
	wire _GEN_2926 = (9'h194 == out_iindex_1 ? _out_T_1122 : _GEN_2925);
	wire _GEN_2927 = (9'h195 == out_iindex_1 ? _out_T_1122 : _GEN_2926);
	wire _GEN_2928 = (9'h196 == out_iindex_1 ? _out_T_1122 : _GEN_2927);
	wire _GEN_2929 = (9'h197 == out_iindex_1 ? _out_T_1122 : _GEN_2928);
	wire _GEN_2930 = (9'h198 == out_iindex_1 ? _out_T_1122 : _GEN_2929);
	wire _GEN_2931 = (9'h199 == out_iindex_1 ? _out_T_1122 : _GEN_2930);
	wire _GEN_2932 = (9'h19a == out_iindex_1 ? _out_T_1122 : _GEN_2931);
	wire _GEN_2933 = (9'h19b == out_iindex_1 ? _out_T_1122 : _GEN_2932);
	wire _GEN_2934 = (9'h19c == out_iindex_1 ? _out_T_1122 : _GEN_2933);
	wire _GEN_2935 = (9'h19d == out_iindex_1 ? _out_T_1122 : _GEN_2934);
	wire _GEN_2936 = (9'h19e == out_iindex_1 ? _out_T_1122 : _GEN_2935);
	wire _GEN_2937 = (9'h19f == out_iindex_1 ? _out_T_1122 : _GEN_2936);
	wire _GEN_2938 = (9'h1a0 == out_iindex_1 ? _out_T_1122 : _GEN_2937);
	wire _GEN_2939 = (9'h1a1 == out_iindex_1 ? _out_T_1122 : _GEN_2938);
	wire _GEN_2940 = (9'h1a2 == out_iindex_1 ? _out_T_1122 : _GEN_2939);
	wire _GEN_2941 = (9'h1a3 == out_iindex_1 ? _out_T_1122 : _GEN_2940);
	wire _GEN_2942 = (9'h1a4 == out_iindex_1 ? _out_T_1122 : _GEN_2941);
	wire _GEN_2943 = (9'h1a5 == out_iindex_1 ? _out_T_1122 : _GEN_2942);
	wire _GEN_2944 = (9'h1a6 == out_iindex_1 ? _out_T_1122 : _GEN_2943);
	wire _GEN_2945 = (9'h1a7 == out_iindex_1 ? _out_T_1122 : _GEN_2944);
	wire _GEN_2946 = (9'h1a8 == out_iindex_1 ? _out_T_1122 : _GEN_2945);
	wire _GEN_2947 = (9'h1a9 == out_iindex_1 ? _out_T_1122 : _GEN_2946);
	wire _GEN_2948 = (9'h1aa == out_iindex_1 ? _out_T_1122 : _GEN_2947);
	wire _GEN_2949 = (9'h1ab == out_iindex_1 ? _out_T_1122 : _GEN_2948);
	wire _GEN_2950 = (9'h1ac == out_iindex_1 ? _out_T_1122 : _GEN_2949);
	wire _GEN_2951 = (9'h1ad == out_iindex_1 ? _out_T_1122 : _GEN_2950);
	wire _GEN_2952 = (9'h1ae == out_iindex_1 ? _out_T_1122 : _GEN_2951);
	wire _GEN_2953 = (9'h1af == out_iindex_1 ? _out_T_1122 : _GEN_2952);
	wire _GEN_2954 = (9'h1b0 == out_iindex_1 ? _out_T_1122 : _GEN_2953);
	wire _GEN_2955 = (9'h1b1 == out_iindex_1 ? _out_T_1122 : _GEN_2954);
	wire _GEN_2956 = (9'h1b2 == out_iindex_1 ? _out_T_1122 : _GEN_2955);
	wire _GEN_2957 = (9'h1b3 == out_iindex_1 ? _out_T_1122 : _GEN_2956);
	wire _GEN_2958 = (9'h1b4 == out_iindex_1 ? _out_T_1122 : _GEN_2957);
	wire _GEN_2959 = (9'h1b5 == out_iindex_1 ? _out_T_1122 : _GEN_2958);
	wire _GEN_2960 = (9'h1b6 == out_iindex_1 ? _out_T_1122 : _GEN_2959);
	wire _GEN_2961 = (9'h1b7 == out_iindex_1 ? _out_T_1122 : _GEN_2960);
	wire _GEN_2962 = (9'h1b8 == out_iindex_1 ? _out_T_1122 : _GEN_2961);
	wire _GEN_2963 = (9'h1b9 == out_iindex_1 ? _out_T_1122 : _GEN_2962);
	wire _GEN_2964 = (9'h1ba == out_iindex_1 ? _out_T_1122 : _GEN_2963);
	wire _GEN_2965 = (9'h1bb == out_iindex_1 ? _out_T_1122 : _GEN_2964);
	wire _GEN_2966 = (9'h1bc == out_iindex_1 ? _out_T_1122 : _GEN_2965);
	wire _GEN_2967 = (9'h1bd == out_iindex_1 ? _out_T_1122 : _GEN_2966);
	wire _GEN_2968 = (9'h1be == out_iindex_1 ? _out_T_1122 : _GEN_2967);
	wire _GEN_2969 = (9'h1bf == out_iindex_1 ? _out_T_1122 : _GEN_2968);
	wire _GEN_2970 = (9'h1c0 == out_iindex_1 ? _out_T_1122 : _GEN_2969);
	wire _GEN_2971 = (9'h1c1 == out_iindex_1 ? _out_T_1122 : _GEN_2970);
	wire _GEN_2972 = (9'h1c2 == out_iindex_1 ? _out_T_1122 : _GEN_2971);
	wire _GEN_2973 = (9'h1c3 == out_iindex_1 ? _out_T_1122 : _GEN_2972);
	wire _GEN_2974 = (9'h1c4 == out_iindex_1 ? _out_T_1122 : _GEN_2973);
	wire _GEN_2975 = (9'h1c5 == out_iindex_1 ? _out_T_1122 : _GEN_2974);
	wire _GEN_2976 = (9'h1c6 == out_iindex_1 ? _out_T_1122 : _GEN_2975);
	wire _GEN_2977 = (9'h1c7 == out_iindex_1 ? _out_T_1122 : _GEN_2976);
	wire _GEN_2978 = (9'h1c8 == out_iindex_1 ? _out_T_1122 : _GEN_2977);
	wire _GEN_2979 = (9'h1c9 == out_iindex_1 ? _out_T_1122 : _GEN_2978);
	wire _GEN_2980 = (9'h1ca == out_iindex_1 ? _out_T_1122 : _GEN_2979);
	wire _GEN_2981 = (9'h1cb == out_iindex_1 ? _out_T_1122 : _GEN_2980);
	wire _GEN_2982 = (9'h1cc == out_iindex_1 ? _out_T_1122 : _GEN_2981);
	wire _GEN_2983 = (9'h1cd == out_iindex_1 ? _out_T_1122 : _GEN_2982);
	wire _GEN_2984 = (9'h1ce == out_iindex_1 ? _out_T_1122 : _GEN_2983);
	wire _GEN_2985 = (9'h1cf == out_iindex_1 ? _out_T_1122 : _GEN_2984);
	wire _GEN_2986 = (9'h1d0 == out_iindex_1 ? _out_T_1122 : _GEN_2985);
	wire _GEN_2987 = (9'h1d1 == out_iindex_1 ? _out_T_1122 : _GEN_2986);
	wire _GEN_2988 = (9'h1d2 == out_iindex_1 ? _out_T_1122 : _GEN_2987);
	wire _GEN_2989 = (9'h1d3 == out_iindex_1 ? _out_T_1122 : _GEN_2988);
	wire _GEN_2990 = (9'h1d4 == out_iindex_1 ? _out_T_1122 : _GEN_2989);
	wire _GEN_2991 = (9'h1d5 == out_iindex_1 ? _out_T_1122 : _GEN_2990);
	wire _GEN_2992 = (9'h1d6 == out_iindex_1 ? _out_T_1122 : _GEN_2991);
	wire _GEN_2993 = (9'h1d7 == out_iindex_1 ? _out_T_1122 : _GEN_2992);
	wire _GEN_2994 = (9'h1d8 == out_iindex_1 ? _out_T_1122 : _GEN_2993);
	wire _GEN_2995 = (9'h1d9 == out_iindex_1 ? _out_T_1122 : _GEN_2994);
	wire _GEN_2996 = (9'h1da == out_iindex_1 ? _out_T_1122 : _GEN_2995);
	wire _GEN_2997 = (9'h1db == out_iindex_1 ? _out_T_1122 : _GEN_2996);
	wire _GEN_2998 = (9'h1dc == out_iindex_1 ? _out_T_1122 : _GEN_2997);
	wire _GEN_2999 = (9'h1dd == out_iindex_1 ? _out_T_1122 : _GEN_2998);
	wire _GEN_3000 = (9'h1de == out_iindex_1 ? _out_T_1122 : _GEN_2999);
	wire _GEN_3001 = (9'h1df == out_iindex_1 ? _out_T_1122 : _GEN_3000);
	wire _GEN_3002 = (9'h1e0 == out_iindex_1 ? _out_T_1122 : _GEN_3001);
	wire _GEN_3003 = (9'h1e1 == out_iindex_1 ? _out_T_1122 : _GEN_3002);
	wire _GEN_3004 = (9'h1e2 == out_iindex_1 ? _out_T_1122 : _GEN_3003);
	wire _GEN_3005 = (9'h1e3 == out_iindex_1 ? _out_T_1122 : _GEN_3004);
	wire _GEN_3006 = (9'h1e4 == out_iindex_1 ? _out_T_1122 : _GEN_3005);
	wire _GEN_3007 = (9'h1e5 == out_iindex_1 ? _out_T_1122 : _GEN_3006);
	wire _GEN_3008 = (9'h1e6 == out_iindex_1 ? _out_T_1122 : _GEN_3007);
	wire _GEN_3009 = (9'h1e7 == out_iindex_1 ? _out_T_1122 : _GEN_3008);
	wire _GEN_3010 = (9'h1e8 == out_iindex_1 ? _out_T_1122 : _GEN_3009);
	wire _GEN_3011 = (9'h1e9 == out_iindex_1 ? _out_T_1122 : _GEN_3010);
	wire _GEN_3012 = (9'h1ea == out_iindex_1 ? _out_T_1122 : _GEN_3011);
	wire _GEN_3013 = (9'h1eb == out_iindex_1 ? _out_T_1122 : _GEN_3012);
	wire _GEN_3014 = (9'h1ec == out_iindex_1 ? _out_T_1122 : _GEN_3013);
	wire _GEN_3015 = (9'h1ed == out_iindex_1 ? _out_T_1122 : _GEN_3014);
	wire _GEN_3016 = (9'h1ee == out_iindex_1 ? _out_T_1122 : _GEN_3015);
	wire _GEN_3017 = (9'h1ef == out_iindex_1 ? _out_T_1122 : _GEN_3016);
	wire _GEN_3018 = (9'h1f0 == out_iindex_1 ? _out_T_1122 : _GEN_3017);
	wire _GEN_3019 = (9'h1f1 == out_iindex_1 ? _out_T_1122 : _GEN_3018);
	wire _GEN_3020 = (9'h1f2 == out_iindex_1 ? _out_T_1122 : _GEN_3019);
	wire _GEN_3021 = (9'h1f3 == out_iindex_1 ? _out_T_1122 : _GEN_3020);
	wire _GEN_3022 = (9'h1f4 == out_iindex_1 ? _out_T_1122 : _GEN_3021);
	wire _GEN_3023 = (9'h1f5 == out_iindex_1 ? _out_T_1122 : _GEN_3022);
	wire _GEN_3024 = (9'h1f6 == out_iindex_1 ? _out_T_1122 : _GEN_3023);
	wire _GEN_3025 = (9'h1f7 == out_iindex_1 ? _out_T_1122 : _GEN_3024);
	wire _GEN_3026 = (9'h1f8 == out_iindex_1 ? _out_T_1122 : _GEN_3025);
	wire _GEN_3027 = (9'h1f9 == out_iindex_1 ? _out_T_1122 : _GEN_3026);
	wire _GEN_3028 = (9'h1fa == out_iindex_1 ? _out_T_1122 : _GEN_3027);
	wire _GEN_3029 = (9'h1fb == out_iindex_1 ? _out_T_1122 : _GEN_3028);
	wire _GEN_3030 = (9'h1fc == out_iindex_1 ? _out_T_1122 : _GEN_3029);
	wire _GEN_3031 = (9'h1fd == out_iindex_1 ? _out_T_1122 : _GEN_3030);
	wire _GEN_3032 = (9'h1fe == out_iindex_1 ? _out_T_1122 : _GEN_3031);
	wire _GEN_3033 = (9'h1ff == out_iindex_1 ? _out_T_1122 : _GEN_3032);
	wire [31:0] _GEN_3035 = (9'h001 == out_iindex_1 ? 32'h0380006f : 32'h00c0006f);
	wire [31:0] _GEN_3036 = (9'h002 == out_iindex_1 ? 32'h0440006f : _GEN_3035);
	wire [31:0] _GEN_3037 = (9'h003 == out_iindex_1 ? 32'h0ff0000f : _GEN_3036);
	wire [31:0] _GEN_3038 = (9'h004 == out_iindex_1 ? 32'h7b241073 : _GEN_3037);
	wire [31:0] _GEN_3039 = (9'h005 == out_iindex_1 ? 32'hf1402473 : _GEN_3038);
	wire [31:0] _GEN_3040 = (9'h006 == out_iindex_1 ? 32'h10802023 : _GEN_3039);
	wire [31:0] _GEN_3041 = (9'h007 == out_iindex_1 ? 32'h40044403 : _GEN_3040);
	wire [31:0] _GEN_3042 = (9'h008 == out_iindex_1 ? 32'h00347413 : _GEN_3041);
	wire [31:0] _GEN_3043 = (9'h009 == out_iindex_1 ? 32'hfe0408e3 : _GEN_3042);
	wire [31:0] _GEN_3044 = (9'h00a == out_iindex_1 ? 32'h00147413 : _GEN_3043);
	wire [31:0] _GEN_3045 = (9'h00b == out_iindex_1 ? 32'h00040863 : _GEN_3044);
	wire [31:0] _GEN_3046 = (9'h00c == out_iindex_1 ? 32'h7b202473 : _GEN_3045);
	wire [31:0] _GEN_3047 = (9'h00d == out_iindex_1 ? 32'h10002223 : _GEN_3046);
	wire [31:0] _GEN_3048 = (9'h00e == out_iindex_1 ? 32'h30000067 : _GEN_3047);
	wire [31:0] _GEN_3049 = (9'h00f == out_iindex_1 ? 32'hf1402473 : _GEN_3048);
	wire [31:0] _GEN_3050 = (9'h010 == out_iindex_1 ? 32'h10802423 : _GEN_3049);
	wire [31:0] _GEN_3051 = (9'h011 == out_iindex_1 ? 32'h7b202473 : _GEN_3050);
	wire [31:0] _GEN_3052 = (9'h012 == out_iindex_1 ? 32'h7b200073 : _GEN_3051);
	wire [31:0] _GEN_3053 = (9'h013 == out_iindex_1 ? 32'h10002623 : _GEN_3052);
	wire [31:0] _GEN_3054 = (9'h014 == out_iindex_1 ? 32'h00100073 : _GEN_3053);
	wire [31:0] _GEN_3055 = (9'h015 == out_iindex_1 ? 32'h00000000 : _GEN_3054);
	wire [31:0] _GEN_3056 = (9'h016 == out_iindex_1 ? 32'h00000000 : _GEN_3055);
	wire [31:0] _GEN_3057 = (9'h017 == out_iindex_1 ? 32'h00000000 : _GEN_3056);
	wire [31:0] _GEN_3058 = (9'h018 == out_iindex_1 ? 32'h00000000 : _GEN_3057);
	wire [31:0] _GEN_3059 = (9'h019 == out_iindex_1 ? 32'h00000000 : _GEN_3058);
	wire [31:0] _GEN_3060 = (9'h01a == out_iindex_1 ? 32'h00000000 : _GEN_3059);
	wire [31:0] _GEN_3061 = (9'h01b == out_iindex_1 ? 32'h00000000 : _GEN_3060);
	wire [31:0] _GEN_3062 = (9'h01c == out_iindex_1 ? 32'h00000000 : _GEN_3061);
	wire [31:0] _GEN_3063 = (9'h01d == out_iindex_1 ? 32'h00000000 : _GEN_3062);
	wire [31:0] _GEN_3064 = (9'h01e == out_iindex_1 ? 32'h00000000 : _GEN_3063);
	wire [31:0] _GEN_3065 = (9'h01f == out_iindex_1 ? 32'h00000000 : _GEN_3064);
	wire [31:0] _GEN_3066 = (9'h020 == out_iindex_1 ? 32'h00000000 : _GEN_3065);
	wire [31:0] _GEN_3067 = (9'h021 == out_iindex_1 ? 32'h00000000 : _GEN_3066);
	wire [31:0] _GEN_3068 = (9'h022 == out_iindex_1 ? 32'h00000000 : _GEN_3067);
	wire [31:0] _GEN_3069 = (9'h023 == out_iindex_1 ? 32'h00000000 : _GEN_3068);
	wire [31:0] _GEN_3070 = (9'h024 == out_iindex_1 ? 32'h00000000 : _GEN_3069);
	wire [31:0] _GEN_3071 = (9'h025 == out_iindex_1 ? 32'h00000000 : _GEN_3070);
	wire [31:0] _GEN_3072 = (9'h026 == out_iindex_1 ? 32'h00000000 : _GEN_3071);
	wire [31:0] _GEN_3073 = (9'h027 == out_iindex_1 ? 32'h00000000 : _GEN_3072);
	wire [31:0] _GEN_3074 = (9'h028 == out_iindex_1 ? 32'h00000000 : _GEN_3073);
	wire [31:0] _GEN_3075 = (9'h029 == out_iindex_1 ? 32'h00000000 : _GEN_3074);
	wire [31:0] _GEN_3076 = (9'h02a == out_iindex_1 ? 32'h00000000 : _GEN_3075);
	wire [31:0] _GEN_3077 = (9'h02b == out_iindex_1 ? 32'h00000000 : _GEN_3076);
	wire [31:0] _GEN_3078 = (9'h02c == out_iindex_1 ? 32'h00000000 : _GEN_3077);
	wire [31:0] _GEN_3079 = (9'h02d == out_iindex_1 ? 32'h00000000 : _GEN_3078);
	wire [31:0] _GEN_3080 = (9'h02e == out_iindex_1 ? 32'h00000000 : _GEN_3079);
	wire [31:0] _GEN_3081 = (9'h02f == out_iindex_1 ? 32'h00000000 : _GEN_3080);
	wire [31:0] _GEN_3082 = (9'h030 == out_iindex_1 ? 32'h00000000 : _GEN_3081);
	wire [31:0] _GEN_3083 = (9'h031 == out_iindex_1 ? 32'h00000000 : _GEN_3082);
	wire [31:0] _GEN_3084 = (9'h032 == out_iindex_1 ? 32'h00000000 : _GEN_3083);
	wire [31:0] _GEN_3085 = (9'h033 == out_iindex_1 ? 32'h00000000 : _GEN_3084);
	wire [31:0] _GEN_3086 = (9'h034 == out_iindex_1 ? 32'h00000000 : _GEN_3085);
	wire [31:0] _GEN_3087 = (9'h035 == out_iindex_1 ? 32'h00000000 : _GEN_3086);
	wire [31:0] _GEN_3088 = (9'h036 == out_iindex_1 ? 32'h00000000 : _GEN_3087);
	wire [31:0] _GEN_3089 = (9'h037 == out_iindex_1 ? 32'h00000000 : _GEN_3088);
	wire [31:0] _GEN_3090 = (9'h038 == out_iindex_1 ? 32'h00000000 : _GEN_3089);
	wire [31:0] _GEN_3091 = (9'h039 == out_iindex_1 ? 32'h00000000 : _GEN_3090);
	wire [31:0] _GEN_3092 = (9'h03a == out_iindex_1 ? 32'h00000000 : _GEN_3091);
	wire [31:0] _GEN_3093 = (9'h03b == out_iindex_1 ? 32'h00000000 : _GEN_3092);
	wire [31:0] _GEN_3094 = (9'h03c == out_iindex_1 ? 32'h00000000 : _GEN_3093);
	wire [31:0] _GEN_3095 = (9'h03d == out_iindex_1 ? 32'h00000000 : _GEN_3094);
	wire [31:0] _GEN_3096 = (9'h03e == out_iindex_1 ? 32'h00000000 : _GEN_3095);
	wire [31:0] _GEN_3097 = (9'h03f == out_iindex_1 ? 32'h00000000 : _GEN_3096);
	wire [31:0] _GEN_3098 = (9'h040 == out_iindex_1 ? 32'h00000000 : _GEN_3097);
	wire [31:0] _GEN_3099 = (9'h041 == out_iindex_1 ? 32'h00000000 : _GEN_3098);
	wire [31:0] _GEN_3100 = (9'h042 == out_iindex_1 ? 32'h00000000 : _GEN_3099);
	wire [31:0] _GEN_3101 = (9'h043 == out_iindex_1 ? 32'h00000000 : _GEN_3100);
	wire [31:0] _GEN_3102 = (9'h044 == out_iindex_1 ? 32'h00000000 : _GEN_3101);
	wire [31:0] _GEN_3103 = (9'h045 == out_iindex_1 ? 32'h00000000 : _GEN_3102);
	wire [31:0] _GEN_3104 = (9'h046 == out_iindex_1 ? 32'h00000000 : _GEN_3103);
	wire [31:0] _GEN_3105 = (9'h047 == out_iindex_1 ? 32'h00000000 : _GEN_3104);
	wire [31:0] _GEN_3106 = (9'h048 == out_iindex_1 ? 32'h00000000 : _GEN_3105);
	wire [31:0] _GEN_3107 = (9'h049 == out_iindex_1 ? 32'h00000000 : _GEN_3106);
	wire [31:0] _GEN_3108 = (9'h04a == out_iindex_1 ? 32'h00000000 : _GEN_3107);
	wire [31:0] _GEN_3109 = (9'h04b == out_iindex_1 ? 32'h00000000 : _GEN_3108);
	wire [31:0] _GEN_3110 = (9'h04c == out_iindex_1 ? 32'h00000000 : _GEN_3109);
	wire [31:0] _GEN_3111 = (9'h04d == out_iindex_1 ? 32'h00000000 : _GEN_3110);
	wire [31:0] _GEN_3112 = (9'h04e == out_iindex_1 ? 32'h00000000 : _GEN_3111);
	wire [31:0] _GEN_3113 = (9'h04f == out_iindex_1 ? 32'h00000000 : _GEN_3112);
	wire [31:0] _GEN_3114 = (9'h050 == out_iindex_1 ? 32'h00000000 : _GEN_3113);
	wire [31:0] _GEN_3115 = (9'h051 == out_iindex_1 ? 32'h00000000 : _GEN_3114);
	wire [31:0] _GEN_3116 = (9'h052 == out_iindex_1 ? 32'h00000000 : _GEN_3115);
	wire [31:0] _GEN_3117 = (9'h053 == out_iindex_1 ? 32'h00000000 : _GEN_3116);
	wire [31:0] _GEN_3118 = (9'h054 == out_iindex_1 ? 32'h00000000 : _GEN_3117);
	wire [31:0] _GEN_3119 = (9'h055 == out_iindex_1 ? 32'h00000000 : _GEN_3118);
	wire [31:0] _GEN_3120 = (9'h056 == out_iindex_1 ? 32'h00000000 : _GEN_3119);
	wire [31:0] _GEN_3121 = (9'h057 == out_iindex_1 ? 32'h00000000 : _GEN_3120);
	wire [31:0] _GEN_3122 = (9'h058 == out_iindex_1 ? 32'h00000000 : _GEN_3121);
	wire [31:0] _GEN_3123 = (9'h059 == out_iindex_1 ? 32'h00000000 : _GEN_3122);
	wire [31:0] _GEN_3124 = (9'h05a == out_iindex_1 ? 32'h00000000 : _GEN_3123);
	wire [31:0] _GEN_3125 = (9'h05b == out_iindex_1 ? 32'h00000000 : _GEN_3124);
	wire [31:0] _GEN_3126 = (9'h05c == out_iindex_1 ? 32'h00000000 : _GEN_3125);
	wire [31:0] _GEN_3127 = (9'h05d == out_iindex_1 ? 32'h00000000 : _GEN_3126);
	wire [31:0] _GEN_3128 = (9'h05e == out_iindex_1 ? 32'h00000000 : _GEN_3127);
	wire [31:0] _GEN_3129 = (9'h05f == out_iindex_1 ? 32'h00000000 : _GEN_3128);
	wire [31:0] _GEN_3130 = (9'h060 == out_iindex_1 ? 32'h00000000 : _GEN_3129);
	wire [31:0] _GEN_3131 = (9'h061 == out_iindex_1 ? 32'h00000000 : _GEN_3130);
	wire [31:0] _GEN_3132 = (9'h062 == out_iindex_1 ? 32'h00000000 : _GEN_3131);
	wire [31:0] _GEN_3133 = (9'h063 == out_iindex_1 ? 32'h00000000 : _GEN_3132);
	wire [31:0] _GEN_3134 = (9'h064 == out_iindex_1 ? 32'h00000000 : _GEN_3133);
	wire [31:0] _GEN_3135 = (9'h065 == out_iindex_1 ? 32'h00000000 : _GEN_3134);
	wire [31:0] _GEN_3136 = (9'h066 == out_iindex_1 ? 32'h00000000 : _GEN_3135);
	wire [31:0] _GEN_3137 = (9'h067 == out_iindex_1 ? 32'h00000000 : _GEN_3136);
	wire [31:0] _GEN_3138 = (9'h068 == out_iindex_1 ? 32'h00000000 : _GEN_3137);
	wire [31:0] _GEN_3139 = (9'h069 == out_iindex_1 ? 32'h00000000 : _GEN_3138);
	wire [31:0] _GEN_3140 = (9'h06a == out_iindex_1 ? 32'h00000000 : _GEN_3139);
	wire [31:0] _GEN_3141 = (9'h06b == out_iindex_1 ? 32'h00000000 : _GEN_3140);
	wire [31:0] _GEN_3142 = (9'h06c == out_iindex_1 ? 32'h00000000 : _GEN_3141);
	wire [31:0] _GEN_3143 = (9'h06d == out_iindex_1 ? 32'h00000000 : _GEN_3142);
	wire [31:0] _GEN_3144 = (9'h06e == out_iindex_1 ? 32'h00000000 : _GEN_3143);
	wire [31:0] _GEN_3145 = (9'h06f == out_iindex_1 ? 32'h00000000 : _GEN_3144);
	wire [31:0] _GEN_3146 = (9'h070 == out_iindex_1 ? 32'h00000000 : _GEN_3145);
	wire [31:0] _GEN_3147 = (9'h071 == out_iindex_1 ? 32'h00000000 : _GEN_3146);
	wire [31:0] _GEN_3148 = (9'h072 == out_iindex_1 ? 32'h00000000 : _GEN_3147);
	wire [31:0] _GEN_3149 = (9'h073 == out_iindex_1 ? 32'h00000000 : _GEN_3148);
	wire [31:0] _GEN_3150 = (9'h074 == out_iindex_1 ? 32'h00000000 : _GEN_3149);
	wire [31:0] _GEN_3151 = (9'h075 == out_iindex_1 ? 32'h00000000 : _GEN_3150);
	wire [31:0] _GEN_3152 = (9'h076 == out_iindex_1 ? 32'h00000000 : _GEN_3151);
	wire [31:0] _GEN_3153 = (9'h077 == out_iindex_1 ? 32'h00000000 : _GEN_3152);
	wire [31:0] _GEN_3154 = (9'h078 == out_iindex_1 ? 32'h00000000 : _GEN_3153);
	wire [31:0] _GEN_3155 = (9'h079 == out_iindex_1 ? 32'h00000000 : _GEN_3154);
	wire [31:0] _GEN_3156 = (9'h07a == out_iindex_1 ? 32'h00000000 : _GEN_3155);
	wire [31:0] _GEN_3157 = (9'h07b == out_iindex_1 ? 32'h00000000 : _GEN_3156);
	wire [31:0] _GEN_3158 = (9'h07c == out_iindex_1 ? 32'h00000000 : _GEN_3157);
	wire [31:0] _GEN_3159 = (9'h07d == out_iindex_1 ? 32'h00000000 : _GEN_3158);
	wire [31:0] _GEN_3160 = (9'h07e == out_iindex_1 ? 32'h00000000 : _GEN_3159);
	wire [31:0] _GEN_3161 = (9'h07f == out_iindex_1 ? 32'h00000000 : _GEN_3160);
	wire [31:0] _GEN_3162 = (9'h080 == out_iindex_1 ? 32'h00000000 : _GEN_3161);
	wire [31:0] _GEN_3163 = (9'h081 == out_iindex_1 ? 32'h00000000 : _GEN_3162);
	wire [31:0] _GEN_3164 = (9'h082 == out_iindex_1 ? 32'h00000000 : _GEN_3163);
	wire [31:0] _GEN_3165 = (9'h083 == out_iindex_1 ? 32'h00000000 : _GEN_3164);
	wire [31:0] _GEN_3166 = (9'h084 == out_iindex_1 ? 32'h00000000 : _GEN_3165);
	wire [31:0] _GEN_3167 = (9'h085 == out_iindex_1 ? 32'h00000000 : _GEN_3166);
	wire [31:0] _GEN_3168 = (9'h086 == out_iindex_1 ? 32'h00000000 : _GEN_3167);
	wire [31:0] _GEN_3169 = (9'h087 == out_iindex_1 ? 32'h00000000 : _GEN_3168);
	wire [31:0] _GEN_3170 = (9'h088 == out_iindex_1 ? 32'h00000000 : _GEN_3169);
	wire [31:0] _GEN_3171 = (9'h089 == out_iindex_1 ? 32'h00000000 : _GEN_3170);
	wire [31:0] _GEN_3172 = (9'h08a == out_iindex_1 ? 32'h00000000 : _GEN_3171);
	wire [31:0] _GEN_3173 = (9'h08b == out_iindex_1 ? 32'h00000000 : _GEN_3172);
	wire [31:0] _GEN_3174 = (9'h08c == out_iindex_1 ? 32'h00000000 : _GEN_3173);
	wire [31:0] _GEN_3175 = (9'h08d == out_iindex_1 ? 32'h00000000 : _GEN_3174);
	wire [31:0] _GEN_3176 = (9'h08e == out_iindex_1 ? 32'h00000000 : _GEN_3175);
	wire [31:0] _GEN_3177 = (9'h08f == out_iindex_1 ? 32'h00000000 : _GEN_3176);
	wire [31:0] _GEN_3178 = (9'h090 == out_iindex_1 ? 32'h00000000 : _GEN_3177);
	wire [31:0] _GEN_3179 = (9'h091 == out_iindex_1 ? 32'h00000000 : _GEN_3178);
	wire [31:0] _GEN_3180 = (9'h092 == out_iindex_1 ? 32'h00000000 : _GEN_3179);
	wire [31:0] _GEN_3181 = (9'h093 == out_iindex_1 ? 32'h00000000 : _GEN_3180);
	wire [31:0] _GEN_3182 = (9'h094 == out_iindex_1 ? 32'h00000000 : _GEN_3181);
	wire [31:0] _GEN_3183 = (9'h095 == out_iindex_1 ? 32'h00000000 : _GEN_3182);
	wire [31:0] _GEN_3184 = (9'h096 == out_iindex_1 ? 32'h00000000 : _GEN_3183);
	wire [31:0] _GEN_3185 = (9'h097 == out_iindex_1 ? 32'h00000000 : _GEN_3184);
	wire [31:0] _GEN_3186 = (9'h098 == out_iindex_1 ? 32'h00000000 : _GEN_3185);
	wire [31:0] _GEN_3187 = (9'h099 == out_iindex_1 ? 32'h00000000 : _GEN_3186);
	wire [31:0] _GEN_3188 = (9'h09a == out_iindex_1 ? 32'h00000000 : _GEN_3187);
	wire [31:0] _GEN_3189 = (9'h09b == out_iindex_1 ? 32'h00000000 : _GEN_3188);
	wire [31:0] _GEN_3190 = (9'h09c == out_iindex_1 ? 32'h00000000 : _GEN_3189);
	wire [31:0] _GEN_3191 = (9'h09d == out_iindex_1 ? 32'h00000000 : _GEN_3190);
	wire [31:0] _GEN_3192 = (9'h09e == out_iindex_1 ? 32'h00000000 : _GEN_3191);
	wire [31:0] _GEN_3193 = (9'h09f == out_iindex_1 ? 32'h00000000 : _GEN_3192);
	wire [31:0] _GEN_3194 = (9'h0a0 == out_iindex_1 ? 32'h00000000 : _GEN_3193);
	wire [31:0] _GEN_3195 = (9'h0a1 == out_iindex_1 ? 32'h00000000 : _GEN_3194);
	wire [31:0] _GEN_3196 = (9'h0a2 == out_iindex_1 ? 32'h00000000 : _GEN_3195);
	wire [31:0] _GEN_3197 = (9'h0a3 == out_iindex_1 ? 32'h00000000 : _GEN_3196);
	wire [31:0] _GEN_3198 = (9'h0a4 == out_iindex_1 ? 32'h00000000 : _GEN_3197);
	wire [31:0] _GEN_3199 = (9'h0a5 == out_iindex_1 ? 32'h00000000 : _GEN_3198);
	wire [31:0] _GEN_3200 = (9'h0a6 == out_iindex_1 ? 32'h00000000 : _GEN_3199);
	wire [31:0] _GEN_3201 = (9'h0a7 == out_iindex_1 ? 32'h00000000 : _GEN_3200);
	wire [31:0] _GEN_3202 = (9'h0a8 == out_iindex_1 ? 32'h00000000 : _GEN_3201);
	wire [31:0] _GEN_3203 = (9'h0a9 == out_iindex_1 ? 32'h00000000 : _GEN_3202);
	wire [31:0] _GEN_3204 = (9'h0aa == out_iindex_1 ? 32'h00000000 : _GEN_3203);
	wire [31:0] _GEN_3205 = (9'h0ab == out_iindex_1 ? 32'h00000000 : _GEN_3204);
	wire [31:0] _GEN_3206 = (9'h0ac == out_iindex_1 ? 32'h00000000 : _GEN_3205);
	wire [31:0] _GEN_3207 = (9'h0ad == out_iindex_1 ? 32'h00000000 : _GEN_3206);
	wire [31:0] _GEN_3208 = (9'h0ae == out_iindex_1 ? 32'h00000000 : _GEN_3207);
	wire [31:0] _GEN_3209 = (9'h0af == out_iindex_1 ? 32'h00000000 : _GEN_3208);
	wire [31:0] _GEN_3210 = (9'h0b0 == out_iindex_1 ? 32'h00000000 : _GEN_3209);
	wire [31:0] _GEN_3211 = (9'h0b1 == out_iindex_1 ? 32'h00000000 : _GEN_3210);
	wire [31:0] _GEN_3212 = (9'h0b2 == out_iindex_1 ? 32'h00000000 : _GEN_3211);
	wire [31:0] _GEN_3213 = (9'h0b3 == out_iindex_1 ? 32'h00000000 : _GEN_3212);
	wire [31:0] _GEN_3214 = (9'h0b4 == out_iindex_1 ? 32'h00000000 : _GEN_3213);
	wire [31:0] _GEN_3215 = (9'h0b5 == out_iindex_1 ? 32'h00000000 : _GEN_3214);
	wire [31:0] _GEN_3216 = (9'h0b6 == out_iindex_1 ? 32'h00000000 : _GEN_3215);
	wire [31:0] _GEN_3217 = (9'h0b7 == out_iindex_1 ? 32'h00000000 : _GEN_3216);
	wire [31:0] _GEN_3218 = (9'h0b8 == out_iindex_1 ? 32'h00000000 : _GEN_3217);
	wire [31:0] _GEN_3219 = (9'h0b9 == out_iindex_1 ? 32'h00000000 : _GEN_3218);
	wire [31:0] _GEN_3220 = (9'h0ba == out_iindex_1 ? 32'h00000000 : _GEN_3219);
	wire [31:0] _GEN_3221 = (9'h0bb == out_iindex_1 ? 32'h00000000 : _GEN_3220);
	wire [31:0] _GEN_3222 = (9'h0bc == out_iindex_1 ? 32'h00000000 : _GEN_3221);
	wire [31:0] _GEN_3223 = (9'h0bd == out_iindex_1 ? 32'h00000000 : _GEN_3222);
	wire [31:0] _GEN_3224 = (9'h0be == out_iindex_1 ? 32'h00000000 : _GEN_3223);
	wire [31:0] _GEN_3225 = (9'h0bf == out_iindex_1 ? 32'h00000000 : _GEN_3224);
	wire [31:0] _GEN_3226 = (9'h0c0 == out_iindex_1 ? 32'h0380006f : _GEN_3225);
	wire [31:0] _GEN_3227 = (9'h0c1 == out_iindex_1 ? 32'h00000000 : _GEN_3226);
	wire [31:0] _GEN_3228 = (9'h0c2 == out_iindex_1 ? 32'h00000000 : _GEN_3227);
	wire [31:0] _GEN_3229 = (9'h0c3 == out_iindex_1 ? 32'h00000000 : _GEN_3228);
	wire [31:0] _GEN_3230 = (9'h0c4 == out_iindex_1 ? 32'h00000000 : _GEN_3229);
	wire [31:0] _GEN_3231 = (9'h0c5 == out_iindex_1 ? 32'h00000000 : _GEN_3230);
	wire [31:0] _GEN_3232 = (9'h0c6 == out_iindex_1 ? 32'h00000000 : _GEN_3231);
	wire [31:0] _GEN_3233 = (9'h0c7 == out_iindex_1 ? 32'h00000000 : _GEN_3232);
	wire [31:0] _GEN_3234 = (9'h0c8 == out_iindex_1 ? 32'h00000000 : _GEN_3233);
	wire [31:0] _GEN_3235 = (9'h0c9 == out_iindex_1 ? 32'h00000000 : _GEN_3234);
	wire [31:0] _GEN_3236 = (9'h0ca == out_iindex_1 ? 32'h00000000 : _GEN_3235);
	wire [31:0] _GEN_3237 = (9'h0cb == out_iindex_1 ? 32'h00000000 : _GEN_3236);
	wire [31:0] _GEN_3238 = (9'h0cc == out_iindex_1 ? 32'h00000000 : _GEN_3237);
	wire [31:0] _GEN_3239 = (9'h0cd == out_iindex_1 ? 32'h00000000 : _GEN_3238);
	wire [31:0] _GEN_3240 = (9'h0ce == out_iindex_1 ? abstractGeneratedMem_0 : _GEN_3239);
	wire [31:0] _GEN_3241 = (9'h0cf == out_iindex_1 ? abstractGeneratedMem_1 : _GEN_3240);
	wire [31:0] _GEN_3242 = (9'h0d0 == out_iindex_1 ? out_prepend_22 : _GEN_3241);
	wire [31:0] _GEN_3243 = (9'h0d1 == out_iindex_1 ? out_prepend_16 : _GEN_3242);
	wire [31:0] _GEN_3244 = (9'h0d2 == out_iindex_1 ? out_prepend_25 : _GEN_3243);
	wire [31:0] _GEN_3245 = (9'h0d3 == out_iindex_1 ? out_prepend_61 : _GEN_3244);
	wire [31:0] _GEN_3246 = (9'h0d4 == out_iindex_1 ? out_prepend_70 : _GEN_3245);
	wire [31:0] _GEN_3247 = (9'h0d5 == out_iindex_1 ? out_prepend_7 : _GEN_3246);
	wire [31:0] _GEN_3248 = (9'h0d6 == out_iindex_1 ? out_prepend_13 : _GEN_3247);
	wire [31:0] _GEN_3249 = (9'h0d7 == out_iindex_1 ? out_prepend_58 : _GEN_3248);
	wire [31:0] _GEN_3250 = (9'h0d8 == out_iindex_1 ? out_prepend_67 : _GEN_3249);
	wire [31:0] _GEN_3251 = (9'h0d9 == out_iindex_1 ? out_prepend_19 : _GEN_3250);
	wire [31:0] _GEN_3252 = (9'h0da == out_iindex_1 ? out_prepend_2 : _GEN_3251);
	wire [31:0] _GEN_3253 = (9'h0db == out_iindex_1 ? out_prepend_64 : _GEN_3252);
	wire [31:0] _GEN_3254 = (9'h0dc == out_iindex_1 ? out_prepend_55 : _GEN_3253);
	wire [31:0] _GEN_3255 = (9'h0dd == out_iindex_1 ? out_prepend_28 : _GEN_3254);
	wire [31:0] _GEN_3256 = (9'h0de == out_iindex_1 ? out_prepend_10 : _GEN_3255);
	wire [31:0] _GEN_3257 = (9'h0df == out_iindex_1 ? out_prepend_76 : _GEN_3256);
	wire [31:0] _GEN_3258 = (9'h0e0 == out_iindex_1 ? out_prepend_73 : _GEN_3257);
	wire [31:0] _GEN_3259 = (9'h0e1 == out_iindex_1 ? 32'h00000000 : _GEN_3258);
	wire [31:0] _GEN_3260 = (9'h0e2 == out_iindex_1 ? 32'h00000000 : _GEN_3259);
	wire [31:0] _GEN_3261 = (9'h0e3 == out_iindex_1 ? 32'h00000000 : _GEN_3260);
	wire [31:0] _GEN_3262 = (9'h0e4 == out_iindex_1 ? 32'h00000000 : _GEN_3261);
	wire [31:0] _GEN_3263 = (9'h0e5 == out_iindex_1 ? 32'h00000000 : _GEN_3262);
	wire [31:0] _GEN_3264 = (9'h0e6 == out_iindex_1 ? 32'h00000000 : _GEN_3263);
	wire [31:0] _GEN_3265 = (9'h0e7 == out_iindex_1 ? 32'h00000000 : _GEN_3264);
	wire [31:0] _GEN_3266 = (9'h0e8 == out_iindex_1 ? 32'h00000000 : _GEN_3265);
	wire [31:0] _GEN_3267 = (9'h0e9 == out_iindex_1 ? 32'h00000000 : _GEN_3266);
	wire [31:0] _GEN_3268 = (9'h0ea == out_iindex_1 ? 32'h00000000 : _GEN_3267);
	wire [31:0] _GEN_3269 = (9'h0eb == out_iindex_1 ? 32'h00000000 : _GEN_3268);
	wire [31:0] _GEN_3270 = (9'h0ec == out_iindex_1 ? 32'h00000000 : _GEN_3269);
	wire [31:0] _GEN_3271 = (9'h0ed == out_iindex_1 ? 32'h00000000 : _GEN_3270);
	wire [31:0] _GEN_3272 = (9'h0ee == out_iindex_1 ? 32'h00000000 : _GEN_3271);
	wire [31:0] _GEN_3273 = (9'h0ef == out_iindex_1 ? 32'h00000000 : _GEN_3272);
	wire [31:0] _GEN_3274 = (9'h0f0 == out_iindex_1 ? 32'h00000000 : _GEN_3273);
	wire [31:0] _GEN_3275 = (9'h0f1 == out_iindex_1 ? 32'h00000000 : _GEN_3274);
	wire [31:0] _GEN_3276 = (9'h0f2 == out_iindex_1 ? 32'h00000000 : _GEN_3275);
	wire [31:0] _GEN_3277 = (9'h0f3 == out_iindex_1 ? 32'h00000000 : _GEN_3276);
	wire [31:0] _GEN_3278 = (9'h0f4 == out_iindex_1 ? 32'h00000000 : _GEN_3277);
	wire [31:0] _GEN_3279 = (9'h0f5 == out_iindex_1 ? 32'h00000000 : _GEN_3278);
	wire [31:0] _GEN_3280 = (9'h0f6 == out_iindex_1 ? 32'h00000000 : _GEN_3279);
	wire [31:0] _GEN_3281 = (9'h0f7 == out_iindex_1 ? 32'h00000000 : _GEN_3280);
	wire [31:0] _GEN_3282 = (9'h0f8 == out_iindex_1 ? 32'h00000000 : _GEN_3281);
	wire [31:0] _GEN_3283 = (9'h0f9 == out_iindex_1 ? 32'h00000000 : _GEN_3282);
	wire [31:0] _GEN_3284 = (9'h0fa == out_iindex_1 ? 32'h00000000 : _GEN_3283);
	wire [31:0] _GEN_3285 = (9'h0fb == out_iindex_1 ? 32'h00000000 : _GEN_3284);
	wire [31:0] _GEN_3286 = (9'h0fc == out_iindex_1 ? 32'h00000000 : _GEN_3285);
	wire [31:0] _GEN_3287 = (9'h0fd == out_iindex_1 ? 32'h00000000 : _GEN_3286);
	wire [31:0] _GEN_3288 = (9'h0fe == out_iindex_1 ? 32'h00000000 : _GEN_3287);
	wire [31:0] _GEN_3289 = (9'h0ff == out_iindex_1 ? 32'h00000000 : _GEN_3288);
	wire [31:0] _GEN_3290 = (9'h100 == out_iindex_1 ? out_prepend_79 : _GEN_3289);
	wire [31:0] _GEN_3291 = (9'h101 == out_iindex_1 ? out_prepend_79 : _GEN_3290);
	wire [31:0] _GEN_3292 = (9'h102 == out_iindex_1 ? out_prepend_79 : _GEN_3291);
	wire [31:0] _GEN_3293 = (9'h103 == out_iindex_1 ? out_prepend_79 : _GEN_3292);
	wire [31:0] _GEN_3294 = (9'h104 == out_iindex_1 ? out_prepend_79 : _GEN_3293);
	wire [31:0] _GEN_3295 = (9'h105 == out_iindex_1 ? out_prepend_79 : _GEN_3294);
	wire [31:0] _GEN_3296 = (9'h106 == out_iindex_1 ? out_prepend_79 : _GEN_3295);
	wire [31:0] _GEN_3297 = (9'h107 == out_iindex_1 ? out_prepend_79 : _GEN_3296);
	wire [31:0] _GEN_3298 = (9'h108 == out_iindex_1 ? out_prepend_79 : _GEN_3297);
	wire [31:0] _GEN_3299 = (9'h109 == out_iindex_1 ? out_prepend_79 : _GEN_3298);
	wire [31:0] _GEN_3300 = (9'h10a == out_iindex_1 ? out_prepend_79 : _GEN_3299);
	wire [31:0] _GEN_3301 = (9'h10b == out_iindex_1 ? out_prepend_79 : _GEN_3300);
	wire [31:0] _GEN_3302 = (9'h10c == out_iindex_1 ? out_prepend_79 : _GEN_3301);
	wire [31:0] _GEN_3303 = (9'h10d == out_iindex_1 ? out_prepend_79 : _GEN_3302);
	wire [31:0] _GEN_3304 = (9'h10e == out_iindex_1 ? out_prepend_79 : _GEN_3303);
	wire [31:0] _GEN_3305 = (9'h10f == out_iindex_1 ? out_prepend_79 : _GEN_3304);
	wire [31:0] _GEN_3306 = (9'h110 == out_iindex_1 ? out_prepend_79 : _GEN_3305);
	wire [31:0] _GEN_3307 = (9'h111 == out_iindex_1 ? out_prepend_79 : _GEN_3306);
	wire [31:0] _GEN_3308 = (9'h112 == out_iindex_1 ? out_prepend_79 : _GEN_3307);
	wire [31:0] _GEN_3309 = (9'h113 == out_iindex_1 ? out_prepend_79 : _GEN_3308);
	wire [31:0] _GEN_3310 = (9'h114 == out_iindex_1 ? out_prepend_79 : _GEN_3309);
	wire [31:0] _GEN_3311 = (9'h115 == out_iindex_1 ? out_prepend_79 : _GEN_3310);
	wire [31:0] _GEN_3312 = (9'h116 == out_iindex_1 ? out_prepend_79 : _GEN_3311);
	wire [31:0] _GEN_3313 = (9'h117 == out_iindex_1 ? out_prepend_79 : _GEN_3312);
	wire [31:0] _GEN_3314 = (9'h118 == out_iindex_1 ? out_prepend_79 : _GEN_3313);
	wire [31:0] _GEN_3315 = (9'h119 == out_iindex_1 ? out_prepend_79 : _GEN_3314);
	wire [31:0] _GEN_3316 = (9'h11a == out_iindex_1 ? out_prepend_79 : _GEN_3315);
	wire [31:0] _GEN_3317 = (9'h11b == out_iindex_1 ? out_prepend_79 : _GEN_3316);
	wire [31:0] _GEN_3318 = (9'h11c == out_iindex_1 ? out_prepend_79 : _GEN_3317);
	wire [31:0] _GEN_3319 = (9'h11d == out_iindex_1 ? out_prepend_79 : _GEN_3318);
	wire [31:0] _GEN_3320 = (9'h11e == out_iindex_1 ? out_prepend_79 : _GEN_3319);
	wire [31:0] _GEN_3321 = (9'h11f == out_iindex_1 ? out_prepend_79 : _GEN_3320);
	wire [31:0] _GEN_3322 = (9'h120 == out_iindex_1 ? out_prepend_79 : _GEN_3321);
	wire [31:0] _GEN_3323 = (9'h121 == out_iindex_1 ? out_prepend_79 : _GEN_3322);
	wire [31:0] _GEN_3324 = (9'h122 == out_iindex_1 ? out_prepend_79 : _GEN_3323);
	wire [31:0] _GEN_3325 = (9'h123 == out_iindex_1 ? out_prepend_79 : _GEN_3324);
	wire [31:0] _GEN_3326 = (9'h124 == out_iindex_1 ? out_prepend_79 : _GEN_3325);
	wire [31:0] _GEN_3327 = (9'h125 == out_iindex_1 ? out_prepend_79 : _GEN_3326);
	wire [31:0] _GEN_3328 = (9'h126 == out_iindex_1 ? out_prepend_79 : _GEN_3327);
	wire [31:0] _GEN_3329 = (9'h127 == out_iindex_1 ? out_prepend_79 : _GEN_3328);
	wire [31:0] _GEN_3330 = (9'h128 == out_iindex_1 ? out_prepend_79 : _GEN_3329);
	wire [31:0] _GEN_3331 = (9'h129 == out_iindex_1 ? out_prepend_79 : _GEN_3330);
	wire [31:0] _GEN_3332 = (9'h12a == out_iindex_1 ? out_prepend_79 : _GEN_3331);
	wire [31:0] _GEN_3333 = (9'h12b == out_iindex_1 ? out_prepend_79 : _GEN_3332);
	wire [31:0] _GEN_3334 = (9'h12c == out_iindex_1 ? out_prepend_79 : _GEN_3333);
	wire [31:0] _GEN_3335 = (9'h12d == out_iindex_1 ? out_prepend_79 : _GEN_3334);
	wire [31:0] _GEN_3336 = (9'h12e == out_iindex_1 ? out_prepend_79 : _GEN_3335);
	wire [31:0] _GEN_3337 = (9'h12f == out_iindex_1 ? out_prepend_79 : _GEN_3336);
	wire [31:0] _GEN_3338 = (9'h130 == out_iindex_1 ? out_prepend_79 : _GEN_3337);
	wire [31:0] _GEN_3339 = (9'h131 == out_iindex_1 ? out_prepend_79 : _GEN_3338);
	wire [31:0] _GEN_3340 = (9'h132 == out_iindex_1 ? out_prepend_79 : _GEN_3339);
	wire [31:0] _GEN_3341 = (9'h133 == out_iindex_1 ? out_prepend_79 : _GEN_3340);
	wire [31:0] _GEN_3342 = (9'h134 == out_iindex_1 ? out_prepend_79 : _GEN_3341);
	wire [31:0] _GEN_3343 = (9'h135 == out_iindex_1 ? out_prepend_79 : _GEN_3342);
	wire [31:0] _GEN_3344 = (9'h136 == out_iindex_1 ? out_prepend_79 : _GEN_3343);
	wire [31:0] _GEN_3345 = (9'h137 == out_iindex_1 ? out_prepend_79 : _GEN_3344);
	wire [31:0] _GEN_3346 = (9'h138 == out_iindex_1 ? out_prepend_79 : _GEN_3345);
	wire [31:0] _GEN_3347 = (9'h139 == out_iindex_1 ? out_prepend_79 : _GEN_3346);
	wire [31:0] _GEN_3348 = (9'h13a == out_iindex_1 ? out_prepend_79 : _GEN_3347);
	wire [31:0] _GEN_3349 = (9'h13b == out_iindex_1 ? out_prepend_79 : _GEN_3348);
	wire [31:0] _GEN_3350 = (9'h13c == out_iindex_1 ? out_prepend_79 : _GEN_3349);
	wire [31:0] _GEN_3351 = (9'h13d == out_iindex_1 ? out_prepend_79 : _GEN_3350);
	wire [31:0] _GEN_3352 = (9'h13e == out_iindex_1 ? out_prepend_79 : _GEN_3351);
	wire [31:0] _GEN_3353 = (9'h13f == out_iindex_1 ? out_prepend_79 : _GEN_3352);
	wire [31:0] _GEN_3354 = (9'h140 == out_iindex_1 ? out_prepend_79 : _GEN_3353);
	wire [31:0] _GEN_3355 = (9'h141 == out_iindex_1 ? out_prepend_79 : _GEN_3354);
	wire [31:0] _GEN_3356 = (9'h142 == out_iindex_1 ? out_prepend_79 : _GEN_3355);
	wire [31:0] _GEN_3357 = (9'h143 == out_iindex_1 ? out_prepend_79 : _GEN_3356);
	wire [31:0] _GEN_3358 = (9'h144 == out_iindex_1 ? out_prepend_79 : _GEN_3357);
	wire [31:0] _GEN_3359 = (9'h145 == out_iindex_1 ? out_prepend_79 : _GEN_3358);
	wire [31:0] _GEN_3360 = (9'h146 == out_iindex_1 ? out_prepend_79 : _GEN_3359);
	wire [31:0] _GEN_3361 = (9'h147 == out_iindex_1 ? out_prepend_79 : _GEN_3360);
	wire [31:0] _GEN_3362 = (9'h148 == out_iindex_1 ? out_prepend_79 : _GEN_3361);
	wire [31:0] _GEN_3363 = (9'h149 == out_iindex_1 ? out_prepend_79 : _GEN_3362);
	wire [31:0] _GEN_3364 = (9'h14a == out_iindex_1 ? out_prepend_79 : _GEN_3363);
	wire [31:0] _GEN_3365 = (9'h14b == out_iindex_1 ? out_prepend_79 : _GEN_3364);
	wire [31:0] _GEN_3366 = (9'h14c == out_iindex_1 ? out_prepend_79 : _GEN_3365);
	wire [31:0] _GEN_3367 = (9'h14d == out_iindex_1 ? out_prepend_79 : _GEN_3366);
	wire [31:0] _GEN_3368 = (9'h14e == out_iindex_1 ? out_prepend_79 : _GEN_3367);
	wire [31:0] _GEN_3369 = (9'h14f == out_iindex_1 ? out_prepend_79 : _GEN_3368);
	wire [31:0] _GEN_3370 = (9'h150 == out_iindex_1 ? out_prepend_79 : _GEN_3369);
	wire [31:0] _GEN_3371 = (9'h151 == out_iindex_1 ? out_prepend_79 : _GEN_3370);
	wire [31:0] _GEN_3372 = (9'h152 == out_iindex_1 ? out_prepend_79 : _GEN_3371);
	wire [31:0] _GEN_3373 = (9'h153 == out_iindex_1 ? out_prepend_79 : _GEN_3372);
	wire [31:0] _GEN_3374 = (9'h154 == out_iindex_1 ? out_prepend_79 : _GEN_3373);
	wire [31:0] _GEN_3375 = (9'h155 == out_iindex_1 ? out_prepend_79 : _GEN_3374);
	wire [31:0] _GEN_3376 = (9'h156 == out_iindex_1 ? out_prepend_79 : _GEN_3375);
	wire [31:0] _GEN_3377 = (9'h157 == out_iindex_1 ? out_prepend_79 : _GEN_3376);
	wire [31:0] _GEN_3378 = (9'h158 == out_iindex_1 ? out_prepend_79 : _GEN_3377);
	wire [31:0] _GEN_3379 = (9'h159 == out_iindex_1 ? out_prepend_79 : _GEN_3378);
	wire [31:0] _GEN_3380 = (9'h15a == out_iindex_1 ? out_prepend_79 : _GEN_3379);
	wire [31:0] _GEN_3381 = (9'h15b == out_iindex_1 ? out_prepend_79 : _GEN_3380);
	wire [31:0] _GEN_3382 = (9'h15c == out_iindex_1 ? out_prepend_79 : _GEN_3381);
	wire [31:0] _GEN_3383 = (9'h15d == out_iindex_1 ? out_prepend_79 : _GEN_3382);
	wire [31:0] _GEN_3384 = (9'h15e == out_iindex_1 ? out_prepend_79 : _GEN_3383);
	wire [31:0] _GEN_3385 = (9'h15f == out_iindex_1 ? out_prepend_79 : _GEN_3384);
	wire [31:0] _GEN_3386 = (9'h160 == out_iindex_1 ? out_prepend_79 : _GEN_3385);
	wire [31:0] _GEN_3387 = (9'h161 == out_iindex_1 ? out_prepend_79 : _GEN_3386);
	wire [31:0] _GEN_3388 = (9'h162 == out_iindex_1 ? out_prepend_79 : _GEN_3387);
	wire [31:0] _GEN_3389 = (9'h163 == out_iindex_1 ? out_prepend_79 : _GEN_3388);
	wire [31:0] _GEN_3390 = (9'h164 == out_iindex_1 ? out_prepend_79 : _GEN_3389);
	wire [31:0] _GEN_3391 = (9'h165 == out_iindex_1 ? out_prepend_79 : _GEN_3390);
	wire [31:0] _GEN_3392 = (9'h166 == out_iindex_1 ? out_prepend_79 : _GEN_3391);
	wire [31:0] _GEN_3393 = (9'h167 == out_iindex_1 ? out_prepend_79 : _GEN_3392);
	wire [31:0] _GEN_3394 = (9'h168 == out_iindex_1 ? out_prepend_79 : _GEN_3393);
	wire [31:0] _GEN_3395 = (9'h169 == out_iindex_1 ? out_prepend_79 : _GEN_3394);
	wire [31:0] _GEN_3396 = (9'h16a == out_iindex_1 ? out_prepend_79 : _GEN_3395);
	wire [31:0] _GEN_3397 = (9'h16b == out_iindex_1 ? out_prepend_79 : _GEN_3396);
	wire [31:0] _GEN_3398 = (9'h16c == out_iindex_1 ? out_prepend_79 : _GEN_3397);
	wire [31:0] _GEN_3399 = (9'h16d == out_iindex_1 ? out_prepend_79 : _GEN_3398);
	wire [31:0] _GEN_3400 = (9'h16e == out_iindex_1 ? out_prepend_79 : _GEN_3399);
	wire [31:0] _GEN_3401 = (9'h16f == out_iindex_1 ? out_prepend_79 : _GEN_3400);
	wire [31:0] _GEN_3402 = (9'h170 == out_iindex_1 ? out_prepend_79 : _GEN_3401);
	wire [31:0] _GEN_3403 = (9'h171 == out_iindex_1 ? out_prepend_79 : _GEN_3402);
	wire [31:0] _GEN_3404 = (9'h172 == out_iindex_1 ? out_prepend_79 : _GEN_3403);
	wire [31:0] _GEN_3405 = (9'h173 == out_iindex_1 ? out_prepend_79 : _GEN_3404);
	wire [31:0] _GEN_3406 = (9'h174 == out_iindex_1 ? out_prepend_79 : _GEN_3405);
	wire [31:0] _GEN_3407 = (9'h175 == out_iindex_1 ? out_prepend_79 : _GEN_3406);
	wire [31:0] _GEN_3408 = (9'h176 == out_iindex_1 ? out_prepend_79 : _GEN_3407);
	wire [31:0] _GEN_3409 = (9'h177 == out_iindex_1 ? out_prepend_79 : _GEN_3408);
	wire [31:0] _GEN_3410 = (9'h178 == out_iindex_1 ? out_prepend_79 : _GEN_3409);
	wire [31:0] _GEN_3411 = (9'h179 == out_iindex_1 ? out_prepend_79 : _GEN_3410);
	wire [31:0] _GEN_3412 = (9'h17a == out_iindex_1 ? out_prepend_79 : _GEN_3411);
	wire [31:0] _GEN_3413 = (9'h17b == out_iindex_1 ? out_prepend_79 : _GEN_3412);
	wire [31:0] _GEN_3414 = (9'h17c == out_iindex_1 ? out_prepend_79 : _GEN_3413);
	wire [31:0] _GEN_3415 = (9'h17d == out_iindex_1 ? out_prepend_79 : _GEN_3414);
	wire [31:0] _GEN_3416 = (9'h17e == out_iindex_1 ? out_prepend_79 : _GEN_3415);
	wire [31:0] _GEN_3417 = (9'h17f == out_iindex_1 ? out_prepend_79 : _GEN_3416);
	wire [31:0] _GEN_3418 = (9'h180 == out_iindex_1 ? out_prepend_79 : _GEN_3417);
	wire [31:0] _GEN_3419 = (9'h181 == out_iindex_1 ? out_prepend_79 : _GEN_3418);
	wire [31:0] _GEN_3420 = (9'h182 == out_iindex_1 ? out_prepend_79 : _GEN_3419);
	wire [31:0] _GEN_3421 = (9'h183 == out_iindex_1 ? out_prepend_79 : _GEN_3420);
	wire [31:0] _GEN_3422 = (9'h184 == out_iindex_1 ? out_prepend_79 : _GEN_3421);
	wire [31:0] _GEN_3423 = (9'h185 == out_iindex_1 ? out_prepend_79 : _GEN_3422);
	wire [31:0] _GEN_3424 = (9'h186 == out_iindex_1 ? out_prepend_79 : _GEN_3423);
	wire [31:0] _GEN_3425 = (9'h187 == out_iindex_1 ? out_prepend_79 : _GEN_3424);
	wire [31:0] _GEN_3426 = (9'h188 == out_iindex_1 ? out_prepend_79 : _GEN_3425);
	wire [31:0] _GEN_3427 = (9'h189 == out_iindex_1 ? out_prepend_79 : _GEN_3426);
	wire [31:0] _GEN_3428 = (9'h18a == out_iindex_1 ? out_prepend_79 : _GEN_3427);
	wire [31:0] _GEN_3429 = (9'h18b == out_iindex_1 ? out_prepend_79 : _GEN_3428);
	wire [31:0] _GEN_3430 = (9'h18c == out_iindex_1 ? out_prepend_79 : _GEN_3429);
	wire [31:0] _GEN_3431 = (9'h18d == out_iindex_1 ? out_prepend_79 : _GEN_3430);
	wire [31:0] _GEN_3432 = (9'h18e == out_iindex_1 ? out_prepend_79 : _GEN_3431);
	wire [31:0] _GEN_3433 = (9'h18f == out_iindex_1 ? out_prepend_79 : _GEN_3432);
	wire [31:0] _GEN_3434 = (9'h190 == out_iindex_1 ? out_prepend_79 : _GEN_3433);
	wire [31:0] _GEN_3435 = (9'h191 == out_iindex_1 ? out_prepend_79 : _GEN_3434);
	wire [31:0] _GEN_3436 = (9'h192 == out_iindex_1 ? out_prepend_79 : _GEN_3435);
	wire [31:0] _GEN_3437 = (9'h193 == out_iindex_1 ? out_prepend_79 : _GEN_3436);
	wire [31:0] _GEN_3438 = (9'h194 == out_iindex_1 ? out_prepend_79 : _GEN_3437);
	wire [31:0] _GEN_3439 = (9'h195 == out_iindex_1 ? out_prepend_79 : _GEN_3438);
	wire [31:0] _GEN_3440 = (9'h196 == out_iindex_1 ? out_prepend_79 : _GEN_3439);
	wire [31:0] _GEN_3441 = (9'h197 == out_iindex_1 ? out_prepend_79 : _GEN_3440);
	wire [31:0] _GEN_3442 = (9'h198 == out_iindex_1 ? out_prepend_79 : _GEN_3441);
	wire [31:0] _GEN_3443 = (9'h199 == out_iindex_1 ? out_prepend_79 : _GEN_3442);
	wire [31:0] _GEN_3444 = (9'h19a == out_iindex_1 ? out_prepend_79 : _GEN_3443);
	wire [31:0] _GEN_3445 = (9'h19b == out_iindex_1 ? out_prepend_79 : _GEN_3444);
	wire [31:0] _GEN_3446 = (9'h19c == out_iindex_1 ? out_prepend_79 : _GEN_3445);
	wire [31:0] _GEN_3447 = (9'h19d == out_iindex_1 ? out_prepend_79 : _GEN_3446);
	wire [31:0] _GEN_3448 = (9'h19e == out_iindex_1 ? out_prepend_79 : _GEN_3447);
	wire [31:0] _GEN_3449 = (9'h19f == out_iindex_1 ? out_prepend_79 : _GEN_3448);
	wire [31:0] _GEN_3450 = (9'h1a0 == out_iindex_1 ? out_prepend_79 : _GEN_3449);
	wire [31:0] _GEN_3451 = (9'h1a1 == out_iindex_1 ? out_prepend_79 : _GEN_3450);
	wire [31:0] _GEN_3452 = (9'h1a2 == out_iindex_1 ? out_prepend_79 : _GEN_3451);
	wire [31:0] _GEN_3453 = (9'h1a3 == out_iindex_1 ? out_prepend_79 : _GEN_3452);
	wire [31:0] _GEN_3454 = (9'h1a4 == out_iindex_1 ? out_prepend_79 : _GEN_3453);
	wire [31:0] _GEN_3455 = (9'h1a5 == out_iindex_1 ? out_prepend_79 : _GEN_3454);
	wire [31:0] _GEN_3456 = (9'h1a6 == out_iindex_1 ? out_prepend_79 : _GEN_3455);
	wire [31:0] _GEN_3457 = (9'h1a7 == out_iindex_1 ? out_prepend_79 : _GEN_3456);
	wire [31:0] _GEN_3458 = (9'h1a8 == out_iindex_1 ? out_prepend_79 : _GEN_3457);
	wire [31:0] _GEN_3459 = (9'h1a9 == out_iindex_1 ? out_prepend_79 : _GEN_3458);
	wire [31:0] _GEN_3460 = (9'h1aa == out_iindex_1 ? out_prepend_79 : _GEN_3459);
	wire [31:0] _GEN_3461 = (9'h1ab == out_iindex_1 ? out_prepend_79 : _GEN_3460);
	wire [31:0] _GEN_3462 = (9'h1ac == out_iindex_1 ? out_prepend_79 : _GEN_3461);
	wire [31:0] _GEN_3463 = (9'h1ad == out_iindex_1 ? out_prepend_79 : _GEN_3462);
	wire [31:0] _GEN_3464 = (9'h1ae == out_iindex_1 ? out_prepend_79 : _GEN_3463);
	wire [31:0] _GEN_3465 = (9'h1af == out_iindex_1 ? out_prepend_79 : _GEN_3464);
	wire [31:0] _GEN_3466 = (9'h1b0 == out_iindex_1 ? out_prepend_79 : _GEN_3465);
	wire [31:0] _GEN_3467 = (9'h1b1 == out_iindex_1 ? out_prepend_79 : _GEN_3466);
	wire [31:0] _GEN_3468 = (9'h1b2 == out_iindex_1 ? out_prepend_79 : _GEN_3467);
	wire [31:0] _GEN_3469 = (9'h1b3 == out_iindex_1 ? out_prepend_79 : _GEN_3468);
	wire [31:0] _GEN_3470 = (9'h1b4 == out_iindex_1 ? out_prepend_79 : _GEN_3469);
	wire [31:0] _GEN_3471 = (9'h1b5 == out_iindex_1 ? out_prepend_79 : _GEN_3470);
	wire [31:0] _GEN_3472 = (9'h1b6 == out_iindex_1 ? out_prepend_79 : _GEN_3471);
	wire [31:0] _GEN_3473 = (9'h1b7 == out_iindex_1 ? out_prepend_79 : _GEN_3472);
	wire [31:0] _GEN_3474 = (9'h1b8 == out_iindex_1 ? out_prepend_79 : _GEN_3473);
	wire [31:0] _GEN_3475 = (9'h1b9 == out_iindex_1 ? out_prepend_79 : _GEN_3474);
	wire [31:0] _GEN_3476 = (9'h1ba == out_iindex_1 ? out_prepend_79 : _GEN_3475);
	wire [31:0] _GEN_3477 = (9'h1bb == out_iindex_1 ? out_prepend_79 : _GEN_3476);
	wire [31:0] _GEN_3478 = (9'h1bc == out_iindex_1 ? out_prepend_79 : _GEN_3477);
	wire [31:0] _GEN_3479 = (9'h1bd == out_iindex_1 ? out_prepend_79 : _GEN_3478);
	wire [31:0] _GEN_3480 = (9'h1be == out_iindex_1 ? out_prepend_79 : _GEN_3479);
	wire [31:0] _GEN_3481 = (9'h1bf == out_iindex_1 ? out_prepend_79 : _GEN_3480);
	wire [31:0] _GEN_3482 = (9'h1c0 == out_iindex_1 ? out_prepend_79 : _GEN_3481);
	wire [31:0] _GEN_3483 = (9'h1c1 == out_iindex_1 ? out_prepend_79 : _GEN_3482);
	wire [31:0] _GEN_3484 = (9'h1c2 == out_iindex_1 ? out_prepend_79 : _GEN_3483);
	wire [31:0] _GEN_3485 = (9'h1c3 == out_iindex_1 ? out_prepend_79 : _GEN_3484);
	wire [31:0] _GEN_3486 = (9'h1c4 == out_iindex_1 ? out_prepend_79 : _GEN_3485);
	wire [31:0] _GEN_3487 = (9'h1c5 == out_iindex_1 ? out_prepend_79 : _GEN_3486);
	wire [31:0] _GEN_3488 = (9'h1c6 == out_iindex_1 ? out_prepend_79 : _GEN_3487);
	wire [31:0] _GEN_3489 = (9'h1c7 == out_iindex_1 ? out_prepend_79 : _GEN_3488);
	wire [31:0] _GEN_3490 = (9'h1c8 == out_iindex_1 ? out_prepend_79 : _GEN_3489);
	wire [31:0] _GEN_3491 = (9'h1c9 == out_iindex_1 ? out_prepend_79 : _GEN_3490);
	wire [31:0] _GEN_3492 = (9'h1ca == out_iindex_1 ? out_prepend_79 : _GEN_3491);
	wire [31:0] _GEN_3493 = (9'h1cb == out_iindex_1 ? out_prepend_79 : _GEN_3492);
	wire [31:0] _GEN_3494 = (9'h1cc == out_iindex_1 ? out_prepend_79 : _GEN_3493);
	wire [31:0] _GEN_3495 = (9'h1cd == out_iindex_1 ? out_prepend_79 : _GEN_3494);
	wire [31:0] _GEN_3496 = (9'h1ce == out_iindex_1 ? out_prepend_79 : _GEN_3495);
	wire [31:0] _GEN_3497 = (9'h1cf == out_iindex_1 ? out_prepend_79 : _GEN_3496);
	wire [31:0] _GEN_3498 = (9'h1d0 == out_iindex_1 ? out_prepend_79 : _GEN_3497);
	wire [31:0] _GEN_3499 = (9'h1d1 == out_iindex_1 ? out_prepend_79 : _GEN_3498);
	wire [31:0] _GEN_3500 = (9'h1d2 == out_iindex_1 ? out_prepend_79 : _GEN_3499);
	wire [31:0] _GEN_3501 = (9'h1d3 == out_iindex_1 ? out_prepend_79 : _GEN_3500);
	wire [31:0] _GEN_3502 = (9'h1d4 == out_iindex_1 ? out_prepend_79 : _GEN_3501);
	wire [31:0] _GEN_3503 = (9'h1d5 == out_iindex_1 ? out_prepend_79 : _GEN_3502);
	wire [31:0] _GEN_3504 = (9'h1d6 == out_iindex_1 ? out_prepend_79 : _GEN_3503);
	wire [31:0] _GEN_3505 = (9'h1d7 == out_iindex_1 ? out_prepend_79 : _GEN_3504);
	wire [31:0] _GEN_3506 = (9'h1d8 == out_iindex_1 ? out_prepend_79 : _GEN_3505);
	wire [31:0] _GEN_3507 = (9'h1d9 == out_iindex_1 ? out_prepend_79 : _GEN_3506);
	wire [31:0] _GEN_3508 = (9'h1da == out_iindex_1 ? out_prepend_79 : _GEN_3507);
	wire [31:0] _GEN_3509 = (9'h1db == out_iindex_1 ? out_prepend_79 : _GEN_3508);
	wire [31:0] _GEN_3510 = (9'h1dc == out_iindex_1 ? out_prepend_79 : _GEN_3509);
	wire [31:0] _GEN_3511 = (9'h1dd == out_iindex_1 ? out_prepend_79 : _GEN_3510);
	wire [31:0] _GEN_3512 = (9'h1de == out_iindex_1 ? out_prepend_79 : _GEN_3511);
	wire [31:0] _GEN_3513 = (9'h1df == out_iindex_1 ? out_prepend_79 : _GEN_3512);
	wire [31:0] _GEN_3514 = (9'h1e0 == out_iindex_1 ? out_prepend_79 : _GEN_3513);
	wire [31:0] _GEN_3515 = (9'h1e1 == out_iindex_1 ? out_prepend_79 : _GEN_3514);
	wire [31:0] _GEN_3516 = (9'h1e2 == out_iindex_1 ? out_prepend_79 : _GEN_3515);
	wire [31:0] _GEN_3517 = (9'h1e3 == out_iindex_1 ? out_prepend_79 : _GEN_3516);
	wire [31:0] _GEN_3518 = (9'h1e4 == out_iindex_1 ? out_prepend_79 : _GEN_3517);
	wire [31:0] _GEN_3519 = (9'h1e5 == out_iindex_1 ? out_prepend_79 : _GEN_3518);
	wire [31:0] _GEN_3520 = (9'h1e6 == out_iindex_1 ? out_prepend_79 : _GEN_3519);
	wire [31:0] _GEN_3521 = (9'h1e7 == out_iindex_1 ? out_prepend_79 : _GEN_3520);
	wire [31:0] _GEN_3522 = (9'h1e8 == out_iindex_1 ? out_prepend_79 : _GEN_3521);
	wire [31:0] _GEN_3523 = (9'h1e9 == out_iindex_1 ? out_prepend_79 : _GEN_3522);
	wire [31:0] _GEN_3524 = (9'h1ea == out_iindex_1 ? out_prepend_79 : _GEN_3523);
	wire [31:0] _GEN_3525 = (9'h1eb == out_iindex_1 ? out_prepend_79 : _GEN_3524);
	wire [31:0] _GEN_3526 = (9'h1ec == out_iindex_1 ? out_prepend_79 : _GEN_3525);
	wire [31:0] _GEN_3527 = (9'h1ed == out_iindex_1 ? out_prepend_79 : _GEN_3526);
	wire [31:0] _GEN_3528 = (9'h1ee == out_iindex_1 ? out_prepend_79 : _GEN_3527);
	wire [31:0] _GEN_3529 = (9'h1ef == out_iindex_1 ? out_prepend_79 : _GEN_3528);
	wire [31:0] _GEN_3530 = (9'h1f0 == out_iindex_1 ? out_prepend_79 : _GEN_3529);
	wire [31:0] _GEN_3531 = (9'h1f1 == out_iindex_1 ? out_prepend_79 : _GEN_3530);
	wire [31:0] _GEN_3532 = (9'h1f2 == out_iindex_1 ? out_prepend_79 : _GEN_3531);
	wire [31:0] _GEN_3533 = (9'h1f3 == out_iindex_1 ? out_prepend_79 : _GEN_3532);
	wire [31:0] _GEN_3534 = (9'h1f4 == out_iindex_1 ? out_prepend_79 : _GEN_3533);
	wire [31:0] _GEN_3535 = (9'h1f5 == out_iindex_1 ? out_prepend_79 : _GEN_3534);
	wire [31:0] _GEN_3536 = (9'h1f6 == out_iindex_1 ? out_prepend_79 : _GEN_3535);
	wire [31:0] _GEN_3537 = (9'h1f7 == out_iindex_1 ? out_prepend_79 : _GEN_3536);
	wire [31:0] _GEN_3538 = (9'h1f8 == out_iindex_1 ? out_prepend_79 : _GEN_3537);
	wire [31:0] _GEN_3539 = (9'h1f9 == out_iindex_1 ? out_prepend_79 : _GEN_3538);
	wire [31:0] _GEN_3540 = (9'h1fa == out_iindex_1 ? out_prepend_79 : _GEN_3539);
	wire [31:0] _GEN_3541 = (9'h1fb == out_iindex_1 ? out_prepend_79 : _GEN_3540);
	wire [31:0] _GEN_3542 = (9'h1fc == out_iindex_1 ? out_prepend_79 : _GEN_3541);
	wire [31:0] _GEN_3543 = (9'h1fd == out_iindex_1 ? out_prepend_79 : _GEN_3542);
	wire [31:0] _GEN_3544 = (9'h1fe == out_iindex_1 ? out_prepend_79 : _GEN_3543);
	wire [31:0] _GEN_3545 = (9'h1ff == out_iindex_1 ? out_prepend_79 : _GEN_3544);
	wire [1:0] _GEN_3627 = (commandRegBadHaltResume ? 2'h0 : 2'h2);
	wire [1:0] _GEN_3633 = (~goReg & out_f_woready_647 ? 2'h0 : ctrlStateReg);
	wire [1:0] _GEN_3634 = (out_f_woready_941 ? 2'h0 : _GEN_3633);
	wire _T_1393 = ctrlStateReg == 2'h3;
	wire _GEN_3894 = _errorBusy_T & ~_T_1383;
	TLMonitor_41 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	TLMonitor_42 monitor_1(
		.clock(monitor_1_clock),
		.reset(monitor_1_reset),
		.io_in_a_ready(monitor_1_io_in_a_ready),
		.io_in_a_valid(monitor_1_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_1_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_1_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_1_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_1_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_1_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_1_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_1_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_1_io_in_d_ready),
		.io_in_d_valid(monitor_1_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_1_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_1_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_1_io_in_d_bits_source)
	);
	AsyncResetSynchronizerShiftReg_w1_d3_i0 hartIsInResetSync_0_debug_hartReset_0(
		.clock(hartIsInResetSync_0_debug_hartReset_0_clock),
		.reset(hartIsInResetSync_0_debug_hartReset_0_reset),
		.io_d(hartIsInResetSync_0_debug_hartReset_0_io_d),
		.io_q(hartIsInResetSync_0_debug_hartReset_0_io_q)
	);
	assign auto_tl_in_a_ready = auto_tl_in_d_ready;
	assign auto_tl_in_d_valid = auto_tl_in_a_valid;
	assign auto_tl_in_d_bits_opcode = {2'd0, in_1_bits_read};
	assign auto_tl_in_d_bits_size = auto_tl_in_a_bits_size;
	assign auto_tl_in_d_bits_source = auto_tl_in_a_bits_source;
	assign auto_tl_in_d_bits_data = (_GEN_3033 ? _GEN_3545 : 32'h00000000);
	assign auto_dmi_in_a_ready = auto_dmi_in_d_ready;
	assign auto_dmi_in_d_valid = auto_dmi_in_a_valid;
	assign auto_dmi_in_d_bits_opcode = {2'd0, in_bits_read};
	assign auto_dmi_in_d_bits_size = auto_dmi_in_a_bits_size;
	assign auto_dmi_in_d_bits_source = auto_dmi_in_a_bits_source;
	assign auto_dmi_in_d_bits_data = (_GEN_296 ? _GEN_328 : 32'h00000000);
	assign io_innerCtrl_ready = 1'h1;
	assign io_hgDebugInt_0 = hrDebugIntReg_0;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_dmi_in_d_ready;
	assign monitor_io_in_a_valid = auto_dmi_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_dmi_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_dmi_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_dmi_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_dmi_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_dmi_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_dmi_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_dmi_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_dmi_in_d_ready;
	assign monitor_io_in_d_valid = auto_dmi_in_a_valid;
	assign monitor_io_in_d_bits_opcode = {2'd0, in_bits_read};
	assign monitor_io_in_d_bits_size = auto_dmi_in_a_bits_size;
	assign monitor_io_in_d_bits_source = auto_dmi_in_a_bits_source;
	assign monitor_1_clock = clock;
	assign monitor_1_reset = reset;
	assign monitor_1_io_in_a_ready = auto_tl_in_d_ready;
	assign monitor_1_io_in_a_valid = auto_tl_in_a_valid;
	assign monitor_1_io_in_a_bits_opcode = auto_tl_in_a_bits_opcode;
	assign monitor_1_io_in_a_bits_param = auto_tl_in_a_bits_param;
	assign monitor_1_io_in_a_bits_size = auto_tl_in_a_bits_size;
	assign monitor_1_io_in_a_bits_source = auto_tl_in_a_bits_source;
	assign monitor_1_io_in_a_bits_address = auto_tl_in_a_bits_address;
	assign monitor_1_io_in_a_bits_mask = auto_tl_in_a_bits_mask;
	assign monitor_1_io_in_a_bits_corrupt = auto_tl_in_a_bits_corrupt;
	assign monitor_1_io_in_d_ready = auto_tl_in_d_ready;
	assign monitor_1_io_in_d_valid = auto_tl_in_a_valid;
	assign monitor_1_io_in_d_bits_opcode = {2'd0, in_1_bits_read};
	assign monitor_1_io_in_d_bits_size = auto_tl_in_a_bits_size;
	assign monitor_1_io_in_d_bits_source = auto_tl_in_a_bits_source;
	assign hartIsInResetSync_0_debug_hartReset_0_clock = clock;
	assign hartIsInResetSync_0_debug_hartReset_0_reset = reset;
	assign hartIsInResetSync_0_debug_hartReset_0_io_d = io_hartIsInReset_0;
	always @(posedge clock) begin
		haltedBitRegs <= _GEN_65[0];
		resumeReqRegs <= _GEN_66[0];
		if (_T_1)
			haveResetBitRegs <= 1'h0;
		else if (_T_4 & io_innerCtrl_bits_ackhavereset)
			haveResetBitRegs <= (haveResetBitRegs & _resumeAcks_T_1) | hartIsInResetSync_0;
		else
			haveResetBitRegs <= haveResetBitRegs | hartIsInResetSync_0;
		if (reset)
			hrmaskReg_0 <= 1'h0;
		else if (~io_dmactive)
			hrmaskReg_0 <= 1'h0;
		else if (_T_4)
			hrmaskReg_0 <= io_innerCtrl_bits_hrmask_0;
		if (_T_1)
			ABSTRACTCSReg_cmderr <= 3'h0;
		else if (errorBusy)
			ABSTRACTCSReg_cmderr <= 3'h1;
		else if (errorException)
			ABSTRACTCSReg_cmderr <= 3'h3;
		else if (errorUnsupported)
			ABSTRACTCSReg_cmderr <= 3'h2;
		else
			ABSTRACTCSReg_cmderr <= _GEN_38;
		if (_T_1)
			ctrlStateReg <= 2'h0;
		else if (ABSTRACTCSWrEnLegal) begin
			if (wrAccessRegisterCommand | regAccessRegisterCommand)
				ctrlStateReg <= 2'h1;
		end
		else if (ctrlStateReg == 2'h1) begin
			if (commandRegIsUnsupported)
				ctrlStateReg <= 2'h0;
			else
				ctrlStateReg <= _GEN_3627;
		end
		else if (ctrlStateReg == 2'h2)
			ctrlStateReg <= _GEN_3634;
		if (_T_1)
			COMMANDRdData_cmdtype <= 8'h00;
		else if (COMMANDWrEn)
			COMMANDRdData_cmdtype <= COMMANDWrData_cmdtype;
		if (_T_1)
			COMMANDRdData_control <= 24'h000000;
		else if (COMMANDWrEn)
			COMMANDRdData_control <= COMMANDWrData_control;
		if (_T_1)
			ABSTRACTAUTOReg_autoexecdata <= 12'h000;
		else if (out_f_woready_4 & ABSTRACTCSWrEnLegal)
			ABSTRACTAUTOReg_autoexecdata <= _ABSTRACTAUTOReg_autoexecdata_T;
		if (_T_1)
			ABSTRACTAUTOReg_autoexecprogbuf <= 16'h0000;
		else if (out_f_woready_6 & ABSTRACTCSWrEnLegal)
			ABSTRACTAUTOReg_autoexecprogbuf <= ABSTRACTAUTOWrData_autoexecprogbuf;
		if (_T_1)
			abstractDataMem_0 <= 8'h00;
		else if (out_f_wivalid_503)
			abstractDataMem_0 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_92 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_92)
				abstractDataMem_0 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			abstractDataMem_1 <= 8'h00;
		else if (out_f_wivalid_504)
			abstractDataMem_1 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_93 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_93)
				abstractDataMem_1 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			abstractDataMem_2 <= 8'h00;
		else if (out_f_wivalid_505)
			abstractDataMem_2 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_94 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_94)
				abstractDataMem_2 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			abstractDataMem_3 <= 8'h00;
		else if (out_f_wivalid_506)
			abstractDataMem_3 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_95 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_95)
				abstractDataMem_3 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_0 <= 8'h00;
		else if (out_f_wivalid_768)
			programBufferMem_0 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_27 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_27)
				programBufferMem_0 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_1 <= 8'h00;
		else if (out_f_wivalid_769)
			programBufferMem_1 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_28 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_28)
				programBufferMem_1 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_2 <= 8'h00;
		else if (out_f_wivalid_770)
			programBufferMem_2 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_29 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_29)
				programBufferMem_2 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_3 <= 8'h00;
		else if (out_f_wivalid_771)
			programBufferMem_3 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_30 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_30)
				programBufferMem_3 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_4 <= 8'h00;
		else if (out_f_wivalid_885)
			programBufferMem_4 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_19 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_19)
				programBufferMem_4 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_5 <= 8'h00;
		else if (out_f_wivalid_886)
			programBufferMem_5 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_20 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_20)
				programBufferMem_5 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_6 <= 8'h00;
		else if (out_f_wivalid_887)
			programBufferMem_6 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_21 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_21)
				programBufferMem_6 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_7 <= 8'h00;
		else if (out_f_wivalid_888)
			programBufferMem_7 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_22 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_22)
				programBufferMem_7 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_8 <= 8'h00;
		else if (out_f_wivalid_1143)
			programBufferMem_8 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_31 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_31)
				programBufferMem_8 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_9 <= 8'h00;
		else if (out_f_wivalid_1144)
			programBufferMem_9 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_32 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_32)
				programBufferMem_9 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_10 <= 8'h00;
		else if (out_f_wivalid_1145)
			programBufferMem_10 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_33 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_33)
				programBufferMem_10 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_11 <= 8'h00;
		else if (out_f_wivalid_1146)
			programBufferMem_11 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_34 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_34)
				programBufferMem_11 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_12 <= 8'h00;
		else if (out_f_wivalid_300)
			programBufferMem_12 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_74 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_74)
				programBufferMem_12 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_13 <= 8'h00;
		else if (out_f_wivalid_301)
			programBufferMem_13 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_75 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_75)
				programBufferMem_13 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_14 <= 8'h00;
		else if (out_f_wivalid_302)
			programBufferMem_14 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_76 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_76)
				programBufferMem_14 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_15 <= 8'h00;
		else if (out_f_wivalid_303)
			programBufferMem_15 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_77 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_77)
				programBufferMem_15 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_16 <= 8'h00;
		else if (out_f_wivalid_567)
			programBufferMem_16 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_87 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_87)
				programBufferMem_16 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_17 <= 8'h00;
		else if (out_f_wivalid_568)
			programBufferMem_17 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_88 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_88)
				programBufferMem_17 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_18 <= 8'h00;
		else if (out_f_wivalid_569)
			programBufferMem_18 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_89 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_89)
				programBufferMem_18 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_19 <= 8'h00;
		else if (out_f_wivalid_570)
			programBufferMem_19 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_90 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_90)
				programBufferMem_19 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_20 <= 8'h00;
		else if (out_f_wivalid_796)
			programBufferMem_20 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_7 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_7)
				programBufferMem_20 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_21 <= 8'h00;
		else if (out_f_wivalid_797)
			programBufferMem_21 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_8 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_8)
				programBufferMem_21 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_22 <= 8'h00;
		else if (out_f_wivalid_798)
			programBufferMem_22 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_9 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_9)
				programBufferMem_22 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_23 <= 8'h00;
		else if (out_f_wivalid_799)
			programBufferMem_23 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_10 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_10)
				programBufferMem_23 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_24 <= 8'h00;
		else if (out_f_wivalid_1091)
			programBufferMem_24 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_15 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_15)
				programBufferMem_24 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_25 <= 8'h00;
		else if (out_f_wivalid_1092)
			programBufferMem_25 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_16 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_16)
				programBufferMem_25 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_26 <= 8'h00;
		else if (out_f_wivalid_1093)
			programBufferMem_26 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_17 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_17)
				programBufferMem_26 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_27 <= 8'h00;
		else if (out_f_wivalid_1094)
			programBufferMem_27 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_18 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_18)
				programBufferMem_27 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_28 <= 8'h00;
		else if (out_f_wivalid_1259)
			programBufferMem_28 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_70 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_70)
				programBufferMem_28 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_29 <= 8'h00;
		else if (out_f_wivalid_1260)
			programBufferMem_29 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_71 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_71)
				programBufferMem_29 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_30 <= 8'h00;
		else if (out_f_wivalid_1261)
			programBufferMem_30 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_72 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_72)
				programBufferMem_30 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_31 <= 8'h00;
		else if (out_f_wivalid_1262)
			programBufferMem_31 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_73 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_73)
				programBufferMem_31 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_32 <= 8'h00;
		else if (out_f_wivalid_276)
			programBufferMem_32 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_82 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_82)
				programBufferMem_32 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_33 <= 8'h00;
		else if (out_f_wivalid_277)
			programBufferMem_33 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_83 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_83)
				programBufferMem_33 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_34 <= 8'h00;
		else if (out_f_wivalid_278)
			programBufferMem_34 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_84 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_84)
				programBufferMem_34 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_35 <= 8'h00;
		else if (out_f_wivalid_279)
			programBufferMem_35 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_85 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_85)
				programBufferMem_35 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_36 <= 8'h00;
		else if (out_f_wivalid_140)
			programBufferMem_36 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_23 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_23)
				programBufferMem_36 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_37 <= 8'h00;
		else if (out_f_wivalid_141)
			programBufferMem_37 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_24 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_24)
				programBufferMem_37 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_38 <= 8'h00;
		else if (out_f_wivalid_142)
			programBufferMem_38 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_25 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_25)
				programBufferMem_38 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_39 <= 8'h00;
		else if (out_f_wivalid_143)
			programBufferMem_39 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_26 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_26)
				programBufferMem_39 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_40 <= 8'h00;
		else if (out_f_wivalid_1018)
			programBufferMem_40 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready & ABSTRACTCSWrEnLegal)
			if (out_f_woready)
				programBufferMem_40 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_41 <= 8'h00;
		else if (out_f_wivalid_1019)
			programBufferMem_41 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_1 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_1)
				programBufferMem_41 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_42 <= 8'h00;
		else if (out_f_wivalid_1020)
			programBufferMem_42 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_2 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_2)
				programBufferMem_42 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_43 <= 8'h00;
		else if (out_f_wivalid_1021)
			programBufferMem_43 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_3 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_3)
				programBufferMem_43 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_44 <= 8'h00;
		else if (out_f_wivalid_724)
			programBufferMem_44 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_78 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_78)
				programBufferMem_44 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_45 <= 8'h00;
		else if (out_f_wivalid_725)
			programBufferMem_45 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_79 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_79)
				programBufferMem_45 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_46 <= 8'h00;
		else if (out_f_wivalid_726)
			programBufferMem_46 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_80 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_80)
				programBufferMem_46 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_47 <= 8'h00;
		else if (out_f_wivalid_727)
			programBufferMem_47 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_81 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_81)
				programBufferMem_47 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_48 <= 8'h00;
		else if (out_f_wivalid_409)
			programBufferMem_48 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_66 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_66)
				programBufferMem_48 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_49 <= 8'h00;
		else if (out_f_wivalid_410)
			programBufferMem_49 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_67 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_67)
				programBufferMem_49 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_50 <= 8'h00;
		else if (out_f_wivalid_411)
			programBufferMem_50 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_68 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_68)
				programBufferMem_50 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_51 <= 8'h00;
		else if (out_f_wivalid_412)
			programBufferMem_51 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_69 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_69)
				programBufferMem_51 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_52 <= 8'h00;
		else if (out_f_wivalid_332)
			programBufferMem_52 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_35 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_35)
				programBufferMem_52 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_53 <= 8'h00;
		else if (out_f_wivalid_333)
			programBufferMem_53 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_36 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_36)
				programBufferMem_53 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_54 <= 8'h00;
		else if (out_f_wivalid_334)
			programBufferMem_54 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_37 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_37)
				programBufferMem_54 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_55 <= 8'h00;
		else if (out_f_wivalid_335)
			programBufferMem_55 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_38 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_38)
				programBufferMem_55 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_56 <= 8'h00;
		else if (out_f_wivalid_1267)
			programBufferMem_56 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_11 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_11)
				programBufferMem_56 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_57 <= 8'h00;
		else if (out_f_wivalid_1268)
			programBufferMem_57 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_12 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_12)
				programBufferMem_57 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_58 <= 8'h00;
		else if (out_f_wivalid_1269)
			programBufferMem_58 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_13 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_13)
				programBufferMem_58 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_59 <= 8'h00;
		else if (out_f_wivalid_1270)
			programBufferMem_59 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_14 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_14)
				programBufferMem_59 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			programBufferMem_60 <= 8'h00;
		else if (out_f_wivalid_833)
			programBufferMem_60 <= auto_tl_in_a_bits_data[7:0];
		else if (out_f_woready_96 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_96)
				programBufferMem_60 <= auto_dmi_in_a_bits_data[7:0];
		if (_T_1)
			programBufferMem_61 <= 8'h00;
		else if (out_f_wivalid_834)
			programBufferMem_61 <= auto_tl_in_a_bits_data[15:8];
		else if (out_f_woready_97 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_97)
				programBufferMem_61 <= auto_dmi_in_a_bits_data[15:8];
		if (_T_1)
			programBufferMem_62 <= 8'h00;
		else if (out_f_wivalid_835)
			programBufferMem_62 <= auto_tl_in_a_bits_data[23:16];
		else if (out_f_woready_98 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_98)
				programBufferMem_62 <= auto_dmi_in_a_bits_data[23:16];
		if (_T_1)
			programBufferMem_63 <= 8'h00;
		else if (out_f_wivalid_836)
			programBufferMem_63 <= auto_tl_in_a_bits_data[31:24];
		else if (out_f_woready_99 & ABSTRACTCSWrEnLegal)
			if (out_f_woready_99)
				programBufferMem_63 <= auto_dmi_in_a_bits_data[31:24];
		if (_T_1)
			goReg <= 1'h0;
		else
			goReg <= _GEN_398;
		if (goAbstract)
			if (accessRegisterCommandReg_transfer) begin
				if (accessRegisterCommandReg_write)
					abstractGeneratedMem_0 <= _abstractGeneratedMem_0_T;
				else
					abstractGeneratedMem_0 <= _abstractGeneratedMem_0_T_1;
			end
			else
				abstractGeneratedMem_0 <= 32'h00000013;
		if (goAbstract)
			if (accessRegisterCommandReg_postexec)
				abstractGeneratedMem_1 <= 32'h00000013;
			else
				abstractGeneratedMem_1 <= 32'h00100073;
	end
	always @(posedge clock or posedge reset)
		if (reset)
			hrDebugIntReg_0 <= 1'h0;
		else if (_T_1)
			hrDebugIntReg_0 <= 1'h0;
		else
			hrDebugIntReg_0 <= _T_13;
endmodule
module ClockCrossingReg_w55 (
	clock,
	io_d,
	io_q,
	io_en
);
	input clock;
	input [54:0] io_d;
	output wire [54:0] io_q;
	input io_en;
	reg [54:0] cdc_reg;
	assign io_q = cdc_reg;
	always @(posedge clock)
		if (io_en)
			cdc_reg <= io_d;
endmodule
module AsyncQueueSink_1 (
	clock,
	reset,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_data,
	io_deq_bits_corrupt,
	io_async_mem_0_opcode,
	io_async_mem_0_address,
	io_async_mem_0_data,
	io_async_ridx,
	io_async_widx,
	io_async_safe_ridx_valid,
	io_async_safe_widx_valid,
	io_async_safe_source_reset_n,
	io_async_safe_sink_reset_n
);
	input clock;
	input reset;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [1:0] io_deq_bits_size;
	output wire io_deq_bits_source;
	output wire [8:0] io_deq_bits_address;
	output wire [3:0] io_deq_bits_mask;
	output wire [31:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	input [2:0] io_async_mem_0_opcode;
	input [8:0] io_async_mem_0_address;
	input [31:0] io_async_mem_0_data;
	output wire io_async_ridx;
	input io_async_widx;
	output wire io_async_safe_ridx_valid;
	input io_async_safe_widx_valid;
	input io_async_safe_source_reset_n;
	output wire io_async_safe_sink_reset_n;
	wire widx_widx_gray_clock;
	wire widx_widx_gray_reset;
	wire widx_widx_gray_io_d;
	wire widx_widx_gray_io_q;
	wire io_deq_bits_deq_bits_reg_clock;
	wire [54:0] io_deq_bits_deq_bits_reg_io_d;
	wire [54:0] io_deq_bits_deq_bits_reg_io_q;
	wire io_deq_bits_deq_bits_reg_io_en;
	wire sink_valid_0_io_in;
	wire sink_valid_0_io_out;
	wire sink_valid_0_clock;
	wire sink_valid_0_reset;
	wire sink_valid_1_io_in;
	wire sink_valid_1_io_out;
	wire sink_valid_1_clock;
	wire sink_valid_1_reset;
	wire source_extend_io_in;
	wire source_extend_io_out;
	wire source_extend_clock;
	wire source_extend_reset;
	wire source_valid_io_in;
	wire source_valid_io_out;
	wire source_valid_clock;
	wire source_valid_reset;
	wire _ridx_T_1 = io_deq_ready & io_deq_valid;
	wire source_ready = source_valid_io_out;
	wire _ridx_T_2 = ~source_ready;
	reg ridx_ridx_bin;
	wire ridx_incremented = (_ridx_T_2 ? 1'h0 : ridx_ridx_bin + _ridx_T_1);
	wire widx = widx_widx_gray_io_q;
	wire [45:0] io_deq_bits_deq_bits_reg_io_d_lo = {io_async_mem_0_address, 4'hf, io_async_mem_0_data, 1'h0};
	wire [8:0] io_deq_bits_deq_bits_reg_io_d_hi = {io_async_mem_0_opcode, 3'h0, 3'h4};
	wire [54:0] _io_deq_bits_WIRE_1 = io_deq_bits_deq_bits_reg_io_q;
	reg valid_reg;
	reg ridx_gray;
	AsyncResetSynchronizerShiftReg_w1_d3_i0 widx_widx_gray(
		.clock(widx_widx_gray_clock),
		.reset(widx_widx_gray_reset),
		.io_d(widx_widx_gray_io_d),
		.io_q(widx_widx_gray_io_q)
	);
	ClockCrossingReg_w55 io_deq_bits_deq_bits_reg(
		.clock(io_deq_bits_deq_bits_reg_clock),
		.io_d(io_deq_bits_deq_bits_reg_io_d),
		.io_q(io_deq_bits_deq_bits_reg_io_q),
		.io_en(io_deq_bits_deq_bits_reg_io_en)
	);
	AsyncValidSync sink_valid_0(
		.io_in(sink_valid_0_io_in),
		.io_out(sink_valid_0_io_out),
		.clock(sink_valid_0_clock),
		.reset(sink_valid_0_reset)
	);
	AsyncValidSync sink_valid_1(
		.io_in(sink_valid_1_io_in),
		.io_out(sink_valid_1_io_out),
		.clock(sink_valid_1_clock),
		.reset(sink_valid_1_reset)
	);
	AsyncValidSync source_extend(
		.io_in(source_extend_io_in),
		.io_out(source_extend_io_out),
		.clock(source_extend_clock),
		.reset(source_extend_reset)
	);
	AsyncValidSync source_valid(
		.io_in(source_valid_io_in),
		.io_out(source_valid_io_out),
		.clock(source_valid_clock),
		.reset(source_valid_reset)
	);
	assign io_deq_valid = valid_reg & source_ready;
	assign io_deq_bits_opcode = _io_deq_bits_WIRE_1[54:52];
	assign io_deq_bits_param = _io_deq_bits_WIRE_1[51:49];
	assign io_deq_bits_size = _io_deq_bits_WIRE_1[48:47];
	assign io_deq_bits_source = _io_deq_bits_WIRE_1[46];
	assign io_deq_bits_address = _io_deq_bits_WIRE_1[45:37];
	assign io_deq_bits_mask = _io_deq_bits_WIRE_1[36:33];
	assign io_deq_bits_data = _io_deq_bits_WIRE_1[32:1];
	assign io_deq_bits_corrupt = _io_deq_bits_WIRE_1[0];
	assign io_async_ridx = ridx_gray;
	assign io_async_safe_ridx_valid = sink_valid_1_io_out;
	assign io_async_safe_sink_reset_n = ~reset;
	assign widx_widx_gray_clock = clock;
	assign widx_widx_gray_reset = reset;
	assign widx_widx_gray_io_d = io_async_widx;
	assign io_deq_bits_deq_bits_reg_clock = clock;
	assign io_deq_bits_deq_bits_reg_io_d = {io_deq_bits_deq_bits_reg_io_d_hi, io_deq_bits_deq_bits_reg_io_d_lo};
	assign io_deq_bits_deq_bits_reg_io_en = source_ready & (ridx_incremented != widx);
	assign sink_valid_0_io_in = 1'h1;
	assign sink_valid_0_clock = clock;
	assign sink_valid_0_reset = reset | ~io_async_safe_source_reset_n;
	assign sink_valid_1_io_in = sink_valid_0_io_out;
	assign sink_valid_1_clock = clock;
	assign sink_valid_1_reset = reset | ~io_async_safe_source_reset_n;
	assign source_extend_io_in = io_async_safe_widx_valid;
	assign source_extend_clock = clock;
	assign source_extend_reset = reset | ~io_async_safe_source_reset_n;
	assign source_valid_io_in = source_extend_io_out;
	assign source_valid_clock = clock;
	assign source_valid_reset = reset;
	always @(posedge clock or posedge reset)
		if (reset)
			ridx_ridx_bin <= 1'h0;
		else if (_ridx_T_2)
			ridx_ridx_bin <= 1'h0;
		else
			ridx_ridx_bin <= ridx_ridx_bin + _ridx_T_1;
	always @(posedge clock or posedge reset)
		if (reset)
			valid_reg <= 1'h0;
		else
			valid_reg <= source_ready & (ridx_incremented != widx);
	always @(posedge clock or posedge reset)
		if (reset)
			ridx_gray <= 1'h0;
		else if (_ridx_T_2)
			ridx_gray <= 1'h0;
		else
			ridx_gray <= ridx_ridx_bin + _ridx_T_1;
endmodule
module AsyncQueueSource_2 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_data,
	io_async_mem_0_opcode,
	io_async_mem_0_size,
	io_async_mem_0_source,
	io_async_mem_0_data,
	io_async_ridx,
	io_async_widx,
	io_async_safe_ridx_valid,
	io_async_safe_widx_valid,
	io_async_safe_source_reset_n,
	io_async_safe_sink_reset_n
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [1:0] io_enq_bits_size;
	input io_enq_bits_source;
	input [31:0] io_enq_bits_data;
	output wire [2:0] io_async_mem_0_opcode;
	output wire [1:0] io_async_mem_0_size;
	output wire io_async_mem_0_source;
	output wire [31:0] io_async_mem_0_data;
	input io_async_ridx;
	output wire io_async_widx;
	input io_async_safe_ridx_valid;
	output wire io_async_safe_widx_valid;
	output wire io_async_safe_source_reset_n;
	input io_async_safe_sink_reset_n;
	wire ridx_ridx_gray_clock;
	wire ridx_ridx_gray_reset;
	wire ridx_ridx_gray_io_d;
	wire ridx_ridx_gray_io_q;
	wire source_valid_0_io_in;
	wire source_valid_0_io_out;
	wire source_valid_0_clock;
	wire source_valid_0_reset;
	wire source_valid_1_io_in;
	wire source_valid_1_io_out;
	wire source_valid_1_clock;
	wire source_valid_1_reset;
	wire sink_extend_io_in;
	wire sink_extend_io_out;
	wire sink_extend_clock;
	wire sink_extend_reset;
	wire sink_valid_io_in;
	wire sink_valid_io_out;
	wire sink_valid_clock;
	wire sink_valid_reset;
	reg [2:0] mem_0_opcode;
	reg [1:0] mem_0_size;
	reg mem_0_source;
	reg [31:0] mem_0_data;
	wire _widx_T_1 = io_enq_ready & io_enq_valid;
	wire sink_ready = sink_valid_io_out;
	wire _widx_T_2 = ~sink_ready;
	reg widx_widx_bin;
	wire widx_incremented = (_widx_T_2 ? 1'h0 : widx_widx_bin + _widx_T_1);
	wire ridx = ridx_ridx_gray_io_q;
	reg ready_reg;
	reg widx_gray;
	AsyncResetSynchronizerShiftReg_w1_d3_i0 ridx_ridx_gray(
		.clock(ridx_ridx_gray_clock),
		.reset(ridx_ridx_gray_reset),
		.io_d(ridx_ridx_gray_io_d),
		.io_q(ridx_ridx_gray_io_q)
	);
	AsyncValidSync source_valid_0(
		.io_in(source_valid_0_io_in),
		.io_out(source_valid_0_io_out),
		.clock(source_valid_0_clock),
		.reset(source_valid_0_reset)
	);
	AsyncValidSync source_valid_1(
		.io_in(source_valid_1_io_in),
		.io_out(source_valid_1_io_out),
		.clock(source_valid_1_clock),
		.reset(source_valid_1_reset)
	);
	AsyncValidSync sink_extend(
		.io_in(sink_extend_io_in),
		.io_out(sink_extend_io_out),
		.clock(sink_extend_clock),
		.reset(sink_extend_reset)
	);
	AsyncValidSync sink_valid(
		.io_in(sink_valid_io_in),
		.io_out(sink_valid_io_out),
		.clock(sink_valid_clock),
		.reset(sink_valid_reset)
	);
	assign io_enq_ready = ready_reg & sink_ready;
	assign io_async_mem_0_opcode = mem_0_opcode;
	assign io_async_mem_0_size = mem_0_size;
	assign io_async_mem_0_source = mem_0_source;
	assign io_async_mem_0_data = mem_0_data;
	assign io_async_widx = widx_gray;
	assign io_async_safe_widx_valid = source_valid_1_io_out;
	assign io_async_safe_source_reset_n = ~reset;
	assign ridx_ridx_gray_clock = clock;
	assign ridx_ridx_gray_reset = reset;
	assign ridx_ridx_gray_io_d = io_async_ridx;
	assign source_valid_0_io_in = 1'h1;
	assign source_valid_0_clock = clock;
	assign source_valid_0_reset = reset | ~io_async_safe_sink_reset_n;
	assign source_valid_1_io_in = source_valid_0_io_out;
	assign source_valid_1_clock = clock;
	assign source_valid_1_reset = reset | ~io_async_safe_sink_reset_n;
	assign sink_extend_io_in = io_async_safe_ridx_valid;
	assign sink_extend_clock = clock;
	assign sink_extend_reset = reset | ~io_async_safe_sink_reset_n;
	assign sink_valid_io_in = sink_extend_io_out;
	assign sink_valid_clock = clock;
	assign sink_valid_reset = reset;
	always @(posedge clock) begin
		if (_widx_T_1)
			mem_0_opcode <= io_enq_bits_opcode;
		if (_widx_T_1)
			mem_0_size <= io_enq_bits_size;
		if (_widx_T_1)
			mem_0_source <= io_enq_bits_source;
		if (_widx_T_1)
			mem_0_data <= io_enq_bits_data;
	end
	always @(posedge clock or posedge reset)
		if (reset)
			widx_widx_bin <= 1'h0;
		else if (_widx_T_2)
			widx_widx_bin <= 1'h0;
		else
			widx_widx_bin <= widx_widx_bin + _widx_T_1;
	always @(posedge clock or posedge reset)
		if (reset)
			ready_reg <= 1'h0;
		else
			ready_reg <= sink_ready & (widx_incremented != (ridx ^ 1'h1));
	always @(posedge clock or posedge reset)
		if (reset)
			widx_gray <= 1'h0;
		else if (_widx_T_2)
			widx_gray <= 1'h0;
		else
			widx_gray <= widx_widx_bin + _widx_T_1;
endmodule
module TLAsyncCrossingSink (
	clock,
	reset,
	auto_in_a_mem_0_opcode,
	auto_in_a_mem_0_address,
	auto_in_a_mem_0_data,
	auto_in_a_ridx,
	auto_in_a_widx,
	auto_in_a_safe_ridx_valid,
	auto_in_a_safe_widx_valid,
	auto_in_a_safe_source_reset_n,
	auto_in_a_safe_sink_reset_n,
	auto_in_d_mem_0_opcode,
	auto_in_d_mem_0_size,
	auto_in_d_mem_0_source,
	auto_in_d_mem_0_data,
	auto_in_d_ridx,
	auto_in_d_widx,
	auto_in_d_safe_ridx_valid,
	auto_in_d_safe_widx_valid,
	auto_in_d_safe_source_reset_n,
	auto_in_d_safe_sink_reset_n,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	input clock;
	input reset;
	input [2:0] auto_in_a_mem_0_opcode;
	input [8:0] auto_in_a_mem_0_address;
	input [31:0] auto_in_a_mem_0_data;
	output wire auto_in_a_ridx;
	input auto_in_a_widx;
	output wire auto_in_a_safe_ridx_valid;
	input auto_in_a_safe_widx_valid;
	input auto_in_a_safe_source_reset_n;
	output wire auto_in_a_safe_sink_reset_n;
	output wire [2:0] auto_in_d_mem_0_opcode;
	output wire [1:0] auto_in_d_mem_0_size;
	output wire auto_in_d_mem_0_source;
	output wire [31:0] auto_in_d_mem_0_data;
	input auto_in_d_ridx;
	output wire auto_in_d_widx;
	input auto_in_d_safe_ridx_valid;
	output wire auto_in_d_safe_widx_valid;
	output wire auto_in_d_safe_source_reset_n;
	input auto_in_d_safe_sink_reset_n;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire auto_out_a_bits_source;
	output wire [8:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_size;
	input auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	wire bundleOut_0_a_sink_clock;
	wire bundleOut_0_a_sink_reset;
	wire bundleOut_0_a_sink_io_deq_ready;
	wire bundleOut_0_a_sink_io_deq_valid;
	wire [2:0] bundleOut_0_a_sink_io_deq_bits_opcode;
	wire [2:0] bundleOut_0_a_sink_io_deq_bits_param;
	wire [1:0] bundleOut_0_a_sink_io_deq_bits_size;
	wire bundleOut_0_a_sink_io_deq_bits_source;
	wire [8:0] bundleOut_0_a_sink_io_deq_bits_address;
	wire [3:0] bundleOut_0_a_sink_io_deq_bits_mask;
	wire [31:0] bundleOut_0_a_sink_io_deq_bits_data;
	wire bundleOut_0_a_sink_io_deq_bits_corrupt;
	wire [2:0] bundleOut_0_a_sink_io_async_mem_0_opcode;
	wire [8:0] bundleOut_0_a_sink_io_async_mem_0_address;
	wire [31:0] bundleOut_0_a_sink_io_async_mem_0_data;
	wire bundleOut_0_a_sink_io_async_ridx;
	wire bundleOut_0_a_sink_io_async_widx;
	wire bundleOut_0_a_sink_io_async_safe_ridx_valid;
	wire bundleOut_0_a_sink_io_async_safe_widx_valid;
	wire bundleOut_0_a_sink_io_async_safe_source_reset_n;
	wire bundleOut_0_a_sink_io_async_safe_sink_reset_n;
	wire bundleIn_0_d_source_clock;
	wire bundleIn_0_d_source_reset;
	wire bundleIn_0_d_source_io_enq_ready;
	wire bundleIn_0_d_source_io_enq_valid;
	wire [2:0] bundleIn_0_d_source_io_enq_bits_opcode;
	wire [1:0] bundleIn_0_d_source_io_enq_bits_size;
	wire bundleIn_0_d_source_io_enq_bits_source;
	wire [31:0] bundleIn_0_d_source_io_enq_bits_data;
	wire [2:0] bundleIn_0_d_source_io_async_mem_0_opcode;
	wire [1:0] bundleIn_0_d_source_io_async_mem_0_size;
	wire bundleIn_0_d_source_io_async_mem_0_source;
	wire [31:0] bundleIn_0_d_source_io_async_mem_0_data;
	wire bundleIn_0_d_source_io_async_ridx;
	wire bundleIn_0_d_source_io_async_widx;
	wire bundleIn_0_d_source_io_async_safe_ridx_valid;
	wire bundleIn_0_d_source_io_async_safe_widx_valid;
	wire bundleIn_0_d_source_io_async_safe_source_reset_n;
	wire bundleIn_0_d_source_io_async_safe_sink_reset_n;
	AsyncQueueSink_1 bundleOut_0_a_sink(
		.clock(bundleOut_0_a_sink_clock),
		.reset(bundleOut_0_a_sink_reset),
		.io_deq_ready(bundleOut_0_a_sink_io_deq_ready),
		.io_deq_valid(bundleOut_0_a_sink_io_deq_valid),
		.io_deq_bits_opcode(bundleOut_0_a_sink_io_deq_bits_opcode),
		.io_deq_bits_param(bundleOut_0_a_sink_io_deq_bits_param),
		.io_deq_bits_size(bundleOut_0_a_sink_io_deq_bits_size),
		.io_deq_bits_source(bundleOut_0_a_sink_io_deq_bits_source),
		.io_deq_bits_address(bundleOut_0_a_sink_io_deq_bits_address),
		.io_deq_bits_mask(bundleOut_0_a_sink_io_deq_bits_mask),
		.io_deq_bits_data(bundleOut_0_a_sink_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleOut_0_a_sink_io_deq_bits_corrupt),
		.io_async_mem_0_opcode(bundleOut_0_a_sink_io_async_mem_0_opcode),
		.io_async_mem_0_address(bundleOut_0_a_sink_io_async_mem_0_address),
		.io_async_mem_0_data(bundleOut_0_a_sink_io_async_mem_0_data),
		.io_async_ridx(bundleOut_0_a_sink_io_async_ridx),
		.io_async_widx(bundleOut_0_a_sink_io_async_widx),
		.io_async_safe_ridx_valid(bundleOut_0_a_sink_io_async_safe_ridx_valid),
		.io_async_safe_widx_valid(bundleOut_0_a_sink_io_async_safe_widx_valid),
		.io_async_safe_source_reset_n(bundleOut_0_a_sink_io_async_safe_source_reset_n),
		.io_async_safe_sink_reset_n(bundleOut_0_a_sink_io_async_safe_sink_reset_n)
	);
	AsyncQueueSource_2 bundleIn_0_d_source(
		.clock(bundleIn_0_d_source_clock),
		.reset(bundleIn_0_d_source_reset),
		.io_enq_ready(bundleIn_0_d_source_io_enq_ready),
		.io_enq_valid(bundleIn_0_d_source_io_enq_valid),
		.io_enq_bits_opcode(bundleIn_0_d_source_io_enq_bits_opcode),
		.io_enq_bits_size(bundleIn_0_d_source_io_enq_bits_size),
		.io_enq_bits_source(bundleIn_0_d_source_io_enq_bits_source),
		.io_enq_bits_data(bundleIn_0_d_source_io_enq_bits_data),
		.io_async_mem_0_opcode(bundleIn_0_d_source_io_async_mem_0_opcode),
		.io_async_mem_0_size(bundleIn_0_d_source_io_async_mem_0_size),
		.io_async_mem_0_source(bundleIn_0_d_source_io_async_mem_0_source),
		.io_async_mem_0_data(bundleIn_0_d_source_io_async_mem_0_data),
		.io_async_ridx(bundleIn_0_d_source_io_async_ridx),
		.io_async_widx(bundleIn_0_d_source_io_async_widx),
		.io_async_safe_ridx_valid(bundleIn_0_d_source_io_async_safe_ridx_valid),
		.io_async_safe_widx_valid(bundleIn_0_d_source_io_async_safe_widx_valid),
		.io_async_safe_source_reset_n(bundleIn_0_d_source_io_async_safe_source_reset_n),
		.io_async_safe_sink_reset_n(bundleIn_0_d_source_io_async_safe_sink_reset_n)
	);
	assign auto_in_a_ridx = bundleOut_0_a_sink_io_async_ridx;
	assign auto_in_a_safe_ridx_valid = bundleOut_0_a_sink_io_async_safe_ridx_valid;
	assign auto_in_a_safe_sink_reset_n = bundleOut_0_a_sink_io_async_safe_sink_reset_n;
	assign auto_in_d_mem_0_opcode = bundleIn_0_d_source_io_async_mem_0_opcode;
	assign auto_in_d_mem_0_size = bundleIn_0_d_source_io_async_mem_0_size;
	assign auto_in_d_mem_0_source = bundleIn_0_d_source_io_async_mem_0_source;
	assign auto_in_d_mem_0_data = bundleIn_0_d_source_io_async_mem_0_data;
	assign auto_in_d_widx = bundleIn_0_d_source_io_async_widx;
	assign auto_in_d_safe_widx_valid = bundleIn_0_d_source_io_async_safe_widx_valid;
	assign auto_in_d_safe_source_reset_n = bundleIn_0_d_source_io_async_safe_source_reset_n;
	assign auto_out_a_valid = bundleOut_0_a_sink_io_deq_valid;
	assign auto_out_a_bits_opcode = bundleOut_0_a_sink_io_deq_bits_opcode;
	assign auto_out_a_bits_param = bundleOut_0_a_sink_io_deq_bits_param;
	assign auto_out_a_bits_size = bundleOut_0_a_sink_io_deq_bits_size;
	assign auto_out_a_bits_source = bundleOut_0_a_sink_io_deq_bits_source;
	assign auto_out_a_bits_address = bundleOut_0_a_sink_io_deq_bits_address;
	assign auto_out_a_bits_mask = bundleOut_0_a_sink_io_deq_bits_mask;
	assign auto_out_a_bits_data = bundleOut_0_a_sink_io_deq_bits_data;
	assign auto_out_a_bits_corrupt = bundleOut_0_a_sink_io_deq_bits_corrupt;
	assign auto_out_d_ready = bundleIn_0_d_source_io_enq_ready;
	assign bundleOut_0_a_sink_clock = clock;
	assign bundleOut_0_a_sink_reset = reset;
	assign bundleOut_0_a_sink_io_deq_ready = auto_out_a_ready;
	assign bundleOut_0_a_sink_io_async_mem_0_opcode = auto_in_a_mem_0_opcode;
	assign bundleOut_0_a_sink_io_async_mem_0_address = auto_in_a_mem_0_address;
	assign bundleOut_0_a_sink_io_async_mem_0_data = auto_in_a_mem_0_data;
	assign bundleOut_0_a_sink_io_async_widx = auto_in_a_widx;
	assign bundleOut_0_a_sink_io_async_safe_widx_valid = auto_in_a_safe_widx_valid;
	assign bundleOut_0_a_sink_io_async_safe_source_reset_n = auto_in_a_safe_source_reset_n;
	assign bundleIn_0_d_source_clock = clock;
	assign bundleIn_0_d_source_reset = reset;
	assign bundleIn_0_d_source_io_enq_valid = auto_out_d_valid;
	assign bundleIn_0_d_source_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign bundleIn_0_d_source_io_enq_bits_size = auto_out_d_bits_size;
	assign bundleIn_0_d_source_io_enq_bits_source = auto_out_d_bits_source;
	assign bundleIn_0_d_source_io_enq_bits_data = auto_out_d_bits_data;
	assign bundleIn_0_d_source_io_async_ridx = auto_in_d_ridx;
	assign bundleIn_0_d_source_io_async_safe_ridx_valid = auto_in_d_safe_ridx_valid;
	assign bundleIn_0_d_source_io_async_safe_sink_reset_n = auto_in_d_safe_sink_reset_n;
endmodule
module ClockCrossingReg_w15 (
	clock,
	io_d,
	io_q,
	io_en
);
	input clock;
	input [14:0] io_d;
	output wire [14:0] io_q;
	input io_en;
	reg [14:0] cdc_reg;
	assign io_q = cdc_reg;
	always @(posedge clock)
		if (io_en)
			cdc_reg <= io_d;
endmodule
module AsyncQueueSink_2 (
	clock,
	reset,
	io_deq_valid,
	io_deq_bits_resumereq,
	io_deq_bits_hartsel,
	io_deq_bits_ackhavereset,
	io_deq_bits_hrmask_0,
	io_async_mem_0_resumereq,
	io_async_mem_0_ackhavereset,
	io_async_mem_0_hrmask_0,
	io_async_ridx,
	io_async_widx,
	io_async_safe_ridx_valid,
	io_async_safe_widx_valid,
	io_async_safe_source_reset_n,
	io_async_safe_sink_reset_n
);
	input clock;
	input reset;
	output wire io_deq_valid;
	output wire io_deq_bits_resumereq;
	output wire [9:0] io_deq_bits_hartsel;
	output wire io_deq_bits_ackhavereset;
	output wire io_deq_bits_hrmask_0;
	input io_async_mem_0_resumereq;
	input io_async_mem_0_ackhavereset;
	input io_async_mem_0_hrmask_0;
	output wire io_async_ridx;
	input io_async_widx;
	output wire io_async_safe_ridx_valid;
	input io_async_safe_widx_valid;
	input io_async_safe_source_reset_n;
	output wire io_async_safe_sink_reset_n;
	wire widx_widx_gray_clock;
	wire widx_widx_gray_reset;
	wire widx_widx_gray_io_d;
	wire widx_widx_gray_io_q;
	wire io_deq_bits_deq_bits_reg_clock;
	wire [14:0] io_deq_bits_deq_bits_reg_io_d;
	wire [14:0] io_deq_bits_deq_bits_reg_io_q;
	wire io_deq_bits_deq_bits_reg_io_en;
	wire sink_valid_0_io_in;
	wire sink_valid_0_io_out;
	wire sink_valid_0_clock;
	wire sink_valid_0_reset;
	wire sink_valid_1_io_in;
	wire sink_valid_1_io_out;
	wire sink_valid_1_clock;
	wire sink_valid_1_reset;
	wire source_extend_io_in;
	wire source_extend_io_out;
	wire source_extend_clock;
	wire source_extend_reset;
	wire source_valid_io_in;
	wire source_valid_io_out;
	wire source_valid_clock;
	wire source_valid_reset;
	wire source_ready = source_valid_io_out;
	wire _ridx_T_2 = ~source_ready;
	reg ridx_ridx_bin;
	wire ridx_incremented = (_ridx_T_2 ? 1'h0 : ridx_ridx_bin + io_deq_valid);
	wire widx = widx_widx_gray_io_q;
	wire [2:0] io_deq_bits_deq_bits_reg_io_d_lo = {2'h0, io_async_mem_0_hrmask_0};
	wire [11:0] io_deq_bits_deq_bits_reg_io_d_hi = {io_async_mem_0_resumereq, 10'h000, io_async_mem_0_ackhavereset};
	wire [14:0] _io_deq_bits_WIRE_1 = io_deq_bits_deq_bits_reg_io_q;
	reg valid_reg;
	reg ridx_gray;
	AsyncResetSynchronizerShiftReg_w1_d3_i0 widx_widx_gray(
		.clock(widx_widx_gray_clock),
		.reset(widx_widx_gray_reset),
		.io_d(widx_widx_gray_io_d),
		.io_q(widx_widx_gray_io_q)
	);
	ClockCrossingReg_w15 io_deq_bits_deq_bits_reg(
		.clock(io_deq_bits_deq_bits_reg_clock),
		.io_d(io_deq_bits_deq_bits_reg_io_d),
		.io_q(io_deq_bits_deq_bits_reg_io_q),
		.io_en(io_deq_bits_deq_bits_reg_io_en)
	);
	AsyncValidSync sink_valid_0(
		.io_in(sink_valid_0_io_in),
		.io_out(sink_valid_0_io_out),
		.clock(sink_valid_0_clock),
		.reset(sink_valid_0_reset)
	);
	AsyncValidSync sink_valid_1(
		.io_in(sink_valid_1_io_in),
		.io_out(sink_valid_1_io_out),
		.clock(sink_valid_1_clock),
		.reset(sink_valid_1_reset)
	);
	AsyncValidSync source_extend(
		.io_in(source_extend_io_in),
		.io_out(source_extend_io_out),
		.clock(source_extend_clock),
		.reset(source_extend_reset)
	);
	AsyncValidSync source_valid(
		.io_in(source_valid_io_in),
		.io_out(source_valid_io_out),
		.clock(source_valid_clock),
		.reset(source_valid_reset)
	);
	assign io_deq_valid = valid_reg & source_ready;
	assign io_deq_bits_resumereq = _io_deq_bits_WIRE_1[14];
	assign io_deq_bits_hartsel = _io_deq_bits_WIRE_1[13:4];
	assign io_deq_bits_ackhavereset = _io_deq_bits_WIRE_1[3];
	assign io_deq_bits_hrmask_0 = _io_deq_bits_WIRE_1[0];
	assign io_async_ridx = ridx_gray;
	assign io_async_safe_ridx_valid = sink_valid_1_io_out;
	assign io_async_safe_sink_reset_n = ~reset;
	assign widx_widx_gray_clock = clock;
	assign widx_widx_gray_reset = reset;
	assign widx_widx_gray_io_d = io_async_widx;
	assign io_deq_bits_deq_bits_reg_clock = clock;
	assign io_deq_bits_deq_bits_reg_io_d = {io_deq_bits_deq_bits_reg_io_d_hi, io_deq_bits_deq_bits_reg_io_d_lo};
	assign io_deq_bits_deq_bits_reg_io_en = source_ready & (ridx_incremented != widx);
	assign sink_valid_0_io_in = 1'h1;
	assign sink_valid_0_clock = clock;
	assign sink_valid_0_reset = reset | ~io_async_safe_source_reset_n;
	assign sink_valid_1_io_in = sink_valid_0_io_out;
	assign sink_valid_1_clock = clock;
	assign sink_valid_1_reset = reset | ~io_async_safe_source_reset_n;
	assign source_extend_io_in = io_async_safe_widx_valid;
	assign source_extend_clock = clock;
	assign source_extend_reset = reset | ~io_async_safe_source_reset_n;
	assign source_valid_io_in = source_extend_io_out;
	assign source_valid_clock = clock;
	assign source_valid_reset = reset;
	always @(posedge clock or posedge reset)
		if (reset)
			ridx_ridx_bin <= 1'h0;
		else if (_ridx_T_2)
			ridx_ridx_bin <= 1'h0;
		else
			ridx_ridx_bin <= ridx_ridx_bin + io_deq_valid;
	always @(posedge clock or posedge reset)
		if (reset)
			valid_reg <= 1'h0;
		else
			valid_reg <= source_ready & (ridx_incremented != widx);
	always @(posedge clock or posedge reset)
		if (reset)
			ridx_gray <= 1'h0;
		else if (_ridx_T_2)
			ridx_gray <= 1'h0;
		else
			ridx_gray <= ridx_ridx_bin + io_deq_valid;
endmodule
module TLDebugModuleInnerAsync (
	auto_dmiXing_in_a_mem_0_opcode,
	auto_dmiXing_in_a_mem_0_address,
	auto_dmiXing_in_a_mem_0_data,
	auto_dmiXing_in_a_ridx,
	auto_dmiXing_in_a_widx,
	auto_dmiXing_in_a_safe_ridx_valid,
	auto_dmiXing_in_a_safe_widx_valid,
	auto_dmiXing_in_a_safe_source_reset_n,
	auto_dmiXing_in_a_safe_sink_reset_n,
	auto_dmiXing_in_d_mem_0_opcode,
	auto_dmiXing_in_d_mem_0_size,
	auto_dmiXing_in_d_mem_0_source,
	auto_dmiXing_in_d_mem_0_data,
	auto_dmiXing_in_d_ridx,
	auto_dmiXing_in_d_widx,
	auto_dmiXing_in_d_safe_ridx_valid,
	auto_dmiXing_in_d_safe_widx_valid,
	auto_dmiXing_in_d_safe_source_reset_n,
	auto_dmiXing_in_d_safe_sink_reset_n,
	auto_dmInner_tl_in_a_ready,
	auto_dmInner_tl_in_a_valid,
	auto_dmInner_tl_in_a_bits_opcode,
	auto_dmInner_tl_in_a_bits_param,
	auto_dmInner_tl_in_a_bits_size,
	auto_dmInner_tl_in_a_bits_source,
	auto_dmInner_tl_in_a_bits_address,
	auto_dmInner_tl_in_a_bits_mask,
	auto_dmInner_tl_in_a_bits_data,
	auto_dmInner_tl_in_a_bits_corrupt,
	auto_dmInner_tl_in_d_ready,
	auto_dmInner_tl_in_d_valid,
	auto_dmInner_tl_in_d_bits_opcode,
	auto_dmInner_tl_in_d_bits_size,
	auto_dmInner_tl_in_d_bits_source,
	auto_dmInner_tl_in_d_bits_data,
	io_debug_clock,
	io_debug_reset,
	io_dmactive,
	io_innerCtrl_mem_0_resumereq,
	io_innerCtrl_mem_0_ackhavereset,
	io_innerCtrl_mem_0_hrmask_0,
	io_innerCtrl_ridx,
	io_innerCtrl_widx,
	io_innerCtrl_safe_ridx_valid,
	io_innerCtrl_safe_widx_valid,
	io_innerCtrl_safe_source_reset_n,
	io_innerCtrl_safe_sink_reset_n,
	io_hgDebugInt_0,
	io_hartIsInReset_0
);
	input [2:0] auto_dmiXing_in_a_mem_0_opcode;
	input [8:0] auto_dmiXing_in_a_mem_0_address;
	input [31:0] auto_dmiXing_in_a_mem_0_data;
	output wire auto_dmiXing_in_a_ridx;
	input auto_dmiXing_in_a_widx;
	output wire auto_dmiXing_in_a_safe_ridx_valid;
	input auto_dmiXing_in_a_safe_widx_valid;
	input auto_dmiXing_in_a_safe_source_reset_n;
	output wire auto_dmiXing_in_a_safe_sink_reset_n;
	output wire [2:0] auto_dmiXing_in_d_mem_0_opcode;
	output wire [1:0] auto_dmiXing_in_d_mem_0_size;
	output wire auto_dmiXing_in_d_mem_0_source;
	output wire [31:0] auto_dmiXing_in_d_mem_0_data;
	input auto_dmiXing_in_d_ridx;
	output wire auto_dmiXing_in_d_widx;
	input auto_dmiXing_in_d_safe_ridx_valid;
	output wire auto_dmiXing_in_d_safe_widx_valid;
	output wire auto_dmiXing_in_d_safe_source_reset_n;
	input auto_dmiXing_in_d_safe_sink_reset_n;
	output wire auto_dmInner_tl_in_a_ready;
	input auto_dmInner_tl_in_a_valid;
	input [2:0] auto_dmInner_tl_in_a_bits_opcode;
	input [2:0] auto_dmInner_tl_in_a_bits_param;
	input [1:0] auto_dmInner_tl_in_a_bits_size;
	input [7:0] auto_dmInner_tl_in_a_bits_source;
	input [11:0] auto_dmInner_tl_in_a_bits_address;
	input [3:0] auto_dmInner_tl_in_a_bits_mask;
	input [31:0] auto_dmInner_tl_in_a_bits_data;
	input auto_dmInner_tl_in_a_bits_corrupt;
	input auto_dmInner_tl_in_d_ready;
	output wire auto_dmInner_tl_in_d_valid;
	output wire [2:0] auto_dmInner_tl_in_d_bits_opcode;
	output wire [1:0] auto_dmInner_tl_in_d_bits_size;
	output wire [7:0] auto_dmInner_tl_in_d_bits_source;
	output wire [31:0] auto_dmInner_tl_in_d_bits_data;
	input io_debug_clock;
	input io_debug_reset;
	input io_dmactive;
	input io_innerCtrl_mem_0_resumereq;
	input io_innerCtrl_mem_0_ackhavereset;
	input io_innerCtrl_mem_0_hrmask_0;
	output wire io_innerCtrl_ridx;
	input io_innerCtrl_widx;
	output wire io_innerCtrl_safe_ridx_valid;
	input io_innerCtrl_safe_widx_valid;
	input io_innerCtrl_safe_source_reset_n;
	output wire io_innerCtrl_safe_sink_reset_n;
	output wire io_hgDebugInt_0;
	input io_hartIsInReset_0;
	wire dmInner_clock;
	wire dmInner_reset;
	wire dmInner_auto_tl_in_a_ready;
	wire dmInner_auto_tl_in_a_valid;
	wire [2:0] dmInner_auto_tl_in_a_bits_opcode;
	wire [2:0] dmInner_auto_tl_in_a_bits_param;
	wire [1:0] dmInner_auto_tl_in_a_bits_size;
	wire [7:0] dmInner_auto_tl_in_a_bits_source;
	wire [11:0] dmInner_auto_tl_in_a_bits_address;
	wire [3:0] dmInner_auto_tl_in_a_bits_mask;
	wire [31:0] dmInner_auto_tl_in_a_bits_data;
	wire dmInner_auto_tl_in_a_bits_corrupt;
	wire dmInner_auto_tl_in_d_ready;
	wire dmInner_auto_tl_in_d_valid;
	wire [2:0] dmInner_auto_tl_in_d_bits_opcode;
	wire [1:0] dmInner_auto_tl_in_d_bits_size;
	wire [7:0] dmInner_auto_tl_in_d_bits_source;
	wire [31:0] dmInner_auto_tl_in_d_bits_data;
	wire dmInner_auto_dmi_in_a_ready;
	wire dmInner_auto_dmi_in_a_valid;
	wire [2:0] dmInner_auto_dmi_in_a_bits_opcode;
	wire [2:0] dmInner_auto_dmi_in_a_bits_param;
	wire [1:0] dmInner_auto_dmi_in_a_bits_size;
	wire dmInner_auto_dmi_in_a_bits_source;
	wire [8:0] dmInner_auto_dmi_in_a_bits_address;
	wire [3:0] dmInner_auto_dmi_in_a_bits_mask;
	wire [31:0] dmInner_auto_dmi_in_a_bits_data;
	wire dmInner_auto_dmi_in_a_bits_corrupt;
	wire dmInner_auto_dmi_in_d_ready;
	wire dmInner_auto_dmi_in_d_valid;
	wire [2:0] dmInner_auto_dmi_in_d_bits_opcode;
	wire [1:0] dmInner_auto_dmi_in_d_bits_size;
	wire dmInner_auto_dmi_in_d_bits_source;
	wire [31:0] dmInner_auto_dmi_in_d_bits_data;
	wire dmInner_io_dmactive;
	wire dmInner_io_innerCtrl_ready;
	wire dmInner_io_innerCtrl_valid;
	wire dmInner_io_innerCtrl_bits_resumereq;
	wire [9:0] dmInner_io_innerCtrl_bits_hartsel;
	wire dmInner_io_innerCtrl_bits_ackhavereset;
	wire dmInner_io_innerCtrl_bits_hrmask_0;
	wire dmInner_io_hgDebugInt_0;
	wire dmInner_io_hartIsInReset_0;
	wire dmiXing_clock;
	wire dmiXing_reset;
	wire [2:0] dmiXing_auto_in_a_mem_0_opcode;
	wire [8:0] dmiXing_auto_in_a_mem_0_address;
	wire [31:0] dmiXing_auto_in_a_mem_0_data;
	wire dmiXing_auto_in_a_ridx;
	wire dmiXing_auto_in_a_widx;
	wire dmiXing_auto_in_a_safe_ridx_valid;
	wire dmiXing_auto_in_a_safe_widx_valid;
	wire dmiXing_auto_in_a_safe_source_reset_n;
	wire dmiXing_auto_in_a_safe_sink_reset_n;
	wire [2:0] dmiXing_auto_in_d_mem_0_opcode;
	wire [1:0] dmiXing_auto_in_d_mem_0_size;
	wire dmiXing_auto_in_d_mem_0_source;
	wire [31:0] dmiXing_auto_in_d_mem_0_data;
	wire dmiXing_auto_in_d_ridx;
	wire dmiXing_auto_in_d_widx;
	wire dmiXing_auto_in_d_safe_ridx_valid;
	wire dmiXing_auto_in_d_safe_widx_valid;
	wire dmiXing_auto_in_d_safe_source_reset_n;
	wire dmiXing_auto_in_d_safe_sink_reset_n;
	wire dmiXing_auto_out_a_ready;
	wire dmiXing_auto_out_a_valid;
	wire [2:0] dmiXing_auto_out_a_bits_opcode;
	wire [2:0] dmiXing_auto_out_a_bits_param;
	wire [1:0] dmiXing_auto_out_a_bits_size;
	wire dmiXing_auto_out_a_bits_source;
	wire [8:0] dmiXing_auto_out_a_bits_address;
	wire [3:0] dmiXing_auto_out_a_bits_mask;
	wire [31:0] dmiXing_auto_out_a_bits_data;
	wire dmiXing_auto_out_a_bits_corrupt;
	wire dmiXing_auto_out_d_ready;
	wire dmiXing_auto_out_d_valid;
	wire [2:0] dmiXing_auto_out_d_bits_opcode;
	wire [1:0] dmiXing_auto_out_d_bits_size;
	wire dmiXing_auto_out_d_bits_source;
	wire [31:0] dmiXing_auto_out_d_bits_data;
	wire dmactive_synced_dmactive_synced_dmactiveSync_clock;
	wire dmactive_synced_dmactive_synced_dmactiveSync_reset;
	wire dmactive_synced_dmactive_synced_dmactiveSync_io_d;
	wire dmactive_synced_dmactive_synced_dmactiveSync_io_q;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_clock;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_reset;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_valid;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_resumereq;
	wire [9:0] dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_hartsel;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_ackhavereset;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_hrmask_0;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_async_mem_0_resumereq;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_async_mem_0_ackhavereset;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_async_mem_0_hrmask_0;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_async_ridx;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_async_widx;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_async_safe_ridx_valid;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_async_safe_widx_valid;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_async_safe_source_reset_n;
	wire dmactive_synced_dmInner_io_innerCtrl_sink_io_async_safe_sink_reset_n;
	TLDebugModuleInner dmInner(
		.clock(dmInner_clock),
		.reset(dmInner_reset),
		.auto_tl_in_a_ready(dmInner_auto_tl_in_a_ready),
		.auto_tl_in_a_valid(dmInner_auto_tl_in_a_valid),
		.auto_tl_in_a_bits_opcode(dmInner_auto_tl_in_a_bits_opcode),
		.auto_tl_in_a_bits_param(dmInner_auto_tl_in_a_bits_param),
		.auto_tl_in_a_bits_size(dmInner_auto_tl_in_a_bits_size),
		.auto_tl_in_a_bits_source(dmInner_auto_tl_in_a_bits_source),
		.auto_tl_in_a_bits_address(dmInner_auto_tl_in_a_bits_address),
		.auto_tl_in_a_bits_mask(dmInner_auto_tl_in_a_bits_mask),
		.auto_tl_in_a_bits_data(dmInner_auto_tl_in_a_bits_data),
		.auto_tl_in_a_bits_corrupt(dmInner_auto_tl_in_a_bits_corrupt),
		.auto_tl_in_d_ready(dmInner_auto_tl_in_d_ready),
		.auto_tl_in_d_valid(dmInner_auto_tl_in_d_valid),
		.auto_tl_in_d_bits_opcode(dmInner_auto_tl_in_d_bits_opcode),
		.auto_tl_in_d_bits_size(dmInner_auto_tl_in_d_bits_size),
		.auto_tl_in_d_bits_source(dmInner_auto_tl_in_d_bits_source),
		.auto_tl_in_d_bits_data(dmInner_auto_tl_in_d_bits_data),
		.auto_dmi_in_a_ready(dmInner_auto_dmi_in_a_ready),
		.auto_dmi_in_a_valid(dmInner_auto_dmi_in_a_valid),
		.auto_dmi_in_a_bits_opcode(dmInner_auto_dmi_in_a_bits_opcode),
		.auto_dmi_in_a_bits_param(dmInner_auto_dmi_in_a_bits_param),
		.auto_dmi_in_a_bits_size(dmInner_auto_dmi_in_a_bits_size),
		.auto_dmi_in_a_bits_source(dmInner_auto_dmi_in_a_bits_source),
		.auto_dmi_in_a_bits_address(dmInner_auto_dmi_in_a_bits_address),
		.auto_dmi_in_a_bits_mask(dmInner_auto_dmi_in_a_bits_mask),
		.auto_dmi_in_a_bits_data(dmInner_auto_dmi_in_a_bits_data),
		.auto_dmi_in_a_bits_corrupt(dmInner_auto_dmi_in_a_bits_corrupt),
		.auto_dmi_in_d_ready(dmInner_auto_dmi_in_d_ready),
		.auto_dmi_in_d_valid(dmInner_auto_dmi_in_d_valid),
		.auto_dmi_in_d_bits_opcode(dmInner_auto_dmi_in_d_bits_opcode),
		.auto_dmi_in_d_bits_size(dmInner_auto_dmi_in_d_bits_size),
		.auto_dmi_in_d_bits_source(dmInner_auto_dmi_in_d_bits_source),
		.auto_dmi_in_d_bits_data(dmInner_auto_dmi_in_d_bits_data),
		.io_dmactive(dmInner_io_dmactive),
		.io_innerCtrl_ready(dmInner_io_innerCtrl_ready),
		.io_innerCtrl_valid(dmInner_io_innerCtrl_valid),
		.io_innerCtrl_bits_resumereq(dmInner_io_innerCtrl_bits_resumereq),
		.io_innerCtrl_bits_hartsel(dmInner_io_innerCtrl_bits_hartsel),
		.io_innerCtrl_bits_ackhavereset(dmInner_io_innerCtrl_bits_ackhavereset),
		.io_innerCtrl_bits_hrmask_0(dmInner_io_innerCtrl_bits_hrmask_0),
		.io_hgDebugInt_0(dmInner_io_hgDebugInt_0),
		.io_hartIsInReset_0(dmInner_io_hartIsInReset_0)
	);
	TLAsyncCrossingSink dmiXing(
		.clock(dmiXing_clock),
		.reset(dmiXing_reset),
		.auto_in_a_mem_0_opcode(dmiXing_auto_in_a_mem_0_opcode),
		.auto_in_a_mem_0_address(dmiXing_auto_in_a_mem_0_address),
		.auto_in_a_mem_0_data(dmiXing_auto_in_a_mem_0_data),
		.auto_in_a_ridx(dmiXing_auto_in_a_ridx),
		.auto_in_a_widx(dmiXing_auto_in_a_widx),
		.auto_in_a_safe_ridx_valid(dmiXing_auto_in_a_safe_ridx_valid),
		.auto_in_a_safe_widx_valid(dmiXing_auto_in_a_safe_widx_valid),
		.auto_in_a_safe_source_reset_n(dmiXing_auto_in_a_safe_source_reset_n),
		.auto_in_a_safe_sink_reset_n(dmiXing_auto_in_a_safe_sink_reset_n),
		.auto_in_d_mem_0_opcode(dmiXing_auto_in_d_mem_0_opcode),
		.auto_in_d_mem_0_size(dmiXing_auto_in_d_mem_0_size),
		.auto_in_d_mem_0_source(dmiXing_auto_in_d_mem_0_source),
		.auto_in_d_mem_0_data(dmiXing_auto_in_d_mem_0_data),
		.auto_in_d_ridx(dmiXing_auto_in_d_ridx),
		.auto_in_d_widx(dmiXing_auto_in_d_widx),
		.auto_in_d_safe_ridx_valid(dmiXing_auto_in_d_safe_ridx_valid),
		.auto_in_d_safe_widx_valid(dmiXing_auto_in_d_safe_widx_valid),
		.auto_in_d_safe_source_reset_n(dmiXing_auto_in_d_safe_source_reset_n),
		.auto_in_d_safe_sink_reset_n(dmiXing_auto_in_d_safe_sink_reset_n),
		.auto_out_a_ready(dmiXing_auto_out_a_ready),
		.auto_out_a_valid(dmiXing_auto_out_a_valid),
		.auto_out_a_bits_opcode(dmiXing_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(dmiXing_auto_out_a_bits_param),
		.auto_out_a_bits_size(dmiXing_auto_out_a_bits_size),
		.auto_out_a_bits_source(dmiXing_auto_out_a_bits_source),
		.auto_out_a_bits_address(dmiXing_auto_out_a_bits_address),
		.auto_out_a_bits_mask(dmiXing_auto_out_a_bits_mask),
		.auto_out_a_bits_data(dmiXing_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(dmiXing_auto_out_a_bits_corrupt),
		.auto_out_d_ready(dmiXing_auto_out_d_ready),
		.auto_out_d_valid(dmiXing_auto_out_d_valid),
		.auto_out_d_bits_opcode(dmiXing_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(dmiXing_auto_out_d_bits_size),
		.auto_out_d_bits_source(dmiXing_auto_out_d_bits_source),
		.auto_out_d_bits_data(dmiXing_auto_out_d_bits_data)
	);
	AsyncResetSynchronizerShiftReg_w1_d3_i0 dmactive_synced_dmactive_synced_dmactiveSync(
		.clock(dmactive_synced_dmactive_synced_dmactiveSync_clock),
		.reset(dmactive_synced_dmactive_synced_dmactiveSync_reset),
		.io_d(dmactive_synced_dmactive_synced_dmactiveSync_io_d),
		.io_q(dmactive_synced_dmactive_synced_dmactiveSync_io_q)
	);
	AsyncQueueSink_2 dmactive_synced_dmInner_io_innerCtrl_sink(
		.clock(dmactive_synced_dmInner_io_innerCtrl_sink_clock),
		.reset(dmactive_synced_dmInner_io_innerCtrl_sink_reset),
		.io_deq_valid(dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_valid),
		.io_deq_bits_resumereq(dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_resumereq),
		.io_deq_bits_hartsel(dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_hartsel),
		.io_deq_bits_ackhavereset(dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_ackhavereset),
		.io_deq_bits_hrmask_0(dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_hrmask_0),
		.io_async_mem_0_resumereq(dmactive_synced_dmInner_io_innerCtrl_sink_io_async_mem_0_resumereq),
		.io_async_mem_0_ackhavereset(dmactive_synced_dmInner_io_innerCtrl_sink_io_async_mem_0_ackhavereset),
		.io_async_mem_0_hrmask_0(dmactive_synced_dmInner_io_innerCtrl_sink_io_async_mem_0_hrmask_0),
		.io_async_ridx(dmactive_synced_dmInner_io_innerCtrl_sink_io_async_ridx),
		.io_async_widx(dmactive_synced_dmInner_io_innerCtrl_sink_io_async_widx),
		.io_async_safe_ridx_valid(dmactive_synced_dmInner_io_innerCtrl_sink_io_async_safe_ridx_valid),
		.io_async_safe_widx_valid(dmactive_synced_dmInner_io_innerCtrl_sink_io_async_safe_widx_valid),
		.io_async_safe_source_reset_n(dmactive_synced_dmInner_io_innerCtrl_sink_io_async_safe_source_reset_n),
		.io_async_safe_sink_reset_n(dmactive_synced_dmInner_io_innerCtrl_sink_io_async_safe_sink_reset_n)
	);
	assign auto_dmiXing_in_a_ridx = dmiXing_auto_in_a_ridx;
	assign auto_dmiXing_in_a_safe_ridx_valid = dmiXing_auto_in_a_safe_ridx_valid;
	assign auto_dmiXing_in_a_safe_sink_reset_n = dmiXing_auto_in_a_safe_sink_reset_n;
	assign auto_dmiXing_in_d_mem_0_opcode = dmiXing_auto_in_d_mem_0_opcode;
	assign auto_dmiXing_in_d_mem_0_size = dmiXing_auto_in_d_mem_0_size;
	assign auto_dmiXing_in_d_mem_0_source = dmiXing_auto_in_d_mem_0_source;
	assign auto_dmiXing_in_d_mem_0_data = dmiXing_auto_in_d_mem_0_data;
	assign auto_dmiXing_in_d_widx = dmiXing_auto_in_d_widx;
	assign auto_dmiXing_in_d_safe_widx_valid = dmiXing_auto_in_d_safe_widx_valid;
	assign auto_dmiXing_in_d_safe_source_reset_n = dmiXing_auto_in_d_safe_source_reset_n;
	assign auto_dmInner_tl_in_a_ready = dmInner_auto_tl_in_a_ready;
	assign auto_dmInner_tl_in_d_valid = dmInner_auto_tl_in_d_valid;
	assign auto_dmInner_tl_in_d_bits_opcode = dmInner_auto_tl_in_d_bits_opcode;
	assign auto_dmInner_tl_in_d_bits_size = dmInner_auto_tl_in_d_bits_size;
	assign auto_dmInner_tl_in_d_bits_source = dmInner_auto_tl_in_d_bits_source;
	assign auto_dmInner_tl_in_d_bits_data = dmInner_auto_tl_in_d_bits_data;
	assign io_innerCtrl_ridx = dmactive_synced_dmInner_io_innerCtrl_sink_io_async_ridx;
	assign io_innerCtrl_safe_ridx_valid = dmactive_synced_dmInner_io_innerCtrl_sink_io_async_safe_ridx_valid;
	assign io_innerCtrl_safe_sink_reset_n = dmactive_synced_dmInner_io_innerCtrl_sink_io_async_safe_sink_reset_n;
	assign io_hgDebugInt_0 = dmInner_io_hgDebugInt_0;
	assign dmInner_clock = io_debug_clock;
	assign dmInner_reset = io_debug_reset;
	assign dmInner_auto_tl_in_a_valid = auto_dmInner_tl_in_a_valid;
	assign dmInner_auto_tl_in_a_bits_opcode = auto_dmInner_tl_in_a_bits_opcode;
	assign dmInner_auto_tl_in_a_bits_param = auto_dmInner_tl_in_a_bits_param;
	assign dmInner_auto_tl_in_a_bits_size = auto_dmInner_tl_in_a_bits_size;
	assign dmInner_auto_tl_in_a_bits_source = auto_dmInner_tl_in_a_bits_source;
	assign dmInner_auto_tl_in_a_bits_address = auto_dmInner_tl_in_a_bits_address;
	assign dmInner_auto_tl_in_a_bits_mask = auto_dmInner_tl_in_a_bits_mask;
	assign dmInner_auto_tl_in_a_bits_data = auto_dmInner_tl_in_a_bits_data;
	assign dmInner_auto_tl_in_a_bits_corrupt = auto_dmInner_tl_in_a_bits_corrupt;
	assign dmInner_auto_tl_in_d_ready = auto_dmInner_tl_in_d_ready;
	assign dmInner_auto_dmi_in_a_valid = dmiXing_auto_out_a_valid;
	assign dmInner_auto_dmi_in_a_bits_opcode = dmiXing_auto_out_a_bits_opcode;
	assign dmInner_auto_dmi_in_a_bits_param = dmiXing_auto_out_a_bits_param;
	assign dmInner_auto_dmi_in_a_bits_size = dmiXing_auto_out_a_bits_size;
	assign dmInner_auto_dmi_in_a_bits_source = dmiXing_auto_out_a_bits_source;
	assign dmInner_auto_dmi_in_a_bits_address = dmiXing_auto_out_a_bits_address;
	assign dmInner_auto_dmi_in_a_bits_mask = dmiXing_auto_out_a_bits_mask;
	assign dmInner_auto_dmi_in_a_bits_data = dmiXing_auto_out_a_bits_data;
	assign dmInner_auto_dmi_in_a_bits_corrupt = dmiXing_auto_out_a_bits_corrupt;
	assign dmInner_auto_dmi_in_d_ready = dmiXing_auto_out_d_ready;
	assign dmInner_io_dmactive = dmactive_synced_dmactive_synced_dmactiveSync_io_q;
	assign dmInner_io_innerCtrl_valid = dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_valid;
	assign dmInner_io_innerCtrl_bits_resumereq = dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_resumereq;
	assign dmInner_io_innerCtrl_bits_hartsel = dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_hartsel;
	assign dmInner_io_innerCtrl_bits_ackhavereset = dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_ackhavereset;
	assign dmInner_io_innerCtrl_bits_hrmask_0 = dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_hrmask_0;
	assign dmInner_io_hartIsInReset_0 = io_hartIsInReset_0;
	assign dmiXing_clock = io_debug_clock;
	assign dmiXing_reset = io_debug_reset;
	assign dmiXing_auto_in_a_mem_0_opcode = auto_dmiXing_in_a_mem_0_opcode;
	assign dmiXing_auto_in_a_mem_0_address = auto_dmiXing_in_a_mem_0_address;
	assign dmiXing_auto_in_a_mem_0_data = auto_dmiXing_in_a_mem_0_data;
	assign dmiXing_auto_in_a_widx = auto_dmiXing_in_a_widx;
	assign dmiXing_auto_in_a_safe_widx_valid = auto_dmiXing_in_a_safe_widx_valid;
	assign dmiXing_auto_in_a_safe_source_reset_n = auto_dmiXing_in_a_safe_source_reset_n;
	assign dmiXing_auto_in_d_ridx = auto_dmiXing_in_d_ridx;
	assign dmiXing_auto_in_d_safe_ridx_valid = auto_dmiXing_in_d_safe_ridx_valid;
	assign dmiXing_auto_in_d_safe_sink_reset_n = auto_dmiXing_in_d_safe_sink_reset_n;
	assign dmiXing_auto_out_a_ready = dmInner_auto_dmi_in_a_ready;
	assign dmiXing_auto_out_d_valid = dmInner_auto_dmi_in_d_valid;
	assign dmiXing_auto_out_d_bits_opcode = dmInner_auto_dmi_in_d_bits_opcode;
	assign dmiXing_auto_out_d_bits_size = dmInner_auto_dmi_in_d_bits_size;
	assign dmiXing_auto_out_d_bits_source = dmInner_auto_dmi_in_d_bits_source;
	assign dmiXing_auto_out_d_bits_data = dmInner_auto_dmi_in_d_bits_data;
	assign dmactive_synced_dmactive_synced_dmactiveSync_clock = io_debug_clock;
	assign dmactive_synced_dmactive_synced_dmactiveSync_reset = io_debug_reset;
	assign dmactive_synced_dmactive_synced_dmactiveSync_io_d = io_dmactive;
	assign dmactive_synced_dmInner_io_innerCtrl_sink_clock = io_debug_clock;
	assign dmactive_synced_dmInner_io_innerCtrl_sink_reset = io_debug_reset;
	assign dmactive_synced_dmInner_io_innerCtrl_sink_io_async_mem_0_resumereq = io_innerCtrl_mem_0_resumereq;
	assign dmactive_synced_dmInner_io_innerCtrl_sink_io_async_mem_0_ackhavereset = io_innerCtrl_mem_0_ackhavereset;
	assign dmactive_synced_dmInner_io_innerCtrl_sink_io_async_mem_0_hrmask_0 = io_innerCtrl_mem_0_hrmask_0;
	assign dmactive_synced_dmInner_io_innerCtrl_sink_io_async_widx = io_innerCtrl_widx;
	assign dmactive_synced_dmInner_io_innerCtrl_sink_io_async_safe_widx_valid = io_innerCtrl_safe_widx_valid;
	assign dmactive_synced_dmInner_io_innerCtrl_sink_io_async_safe_source_reset_n = io_innerCtrl_safe_source_reset_n;
endmodule
module TLDebugModule (
	auto_dmInner_dmInner_tl_in_a_ready,
	auto_dmInner_dmInner_tl_in_a_valid,
	auto_dmInner_dmInner_tl_in_a_bits_opcode,
	auto_dmInner_dmInner_tl_in_a_bits_param,
	auto_dmInner_dmInner_tl_in_a_bits_size,
	auto_dmInner_dmInner_tl_in_a_bits_source,
	auto_dmInner_dmInner_tl_in_a_bits_address,
	auto_dmInner_dmInner_tl_in_a_bits_mask,
	auto_dmInner_dmInner_tl_in_a_bits_data,
	auto_dmInner_dmInner_tl_in_a_bits_corrupt,
	auto_dmInner_dmInner_tl_in_d_ready,
	auto_dmInner_dmInner_tl_in_d_valid,
	auto_dmInner_dmInner_tl_in_d_bits_opcode,
	auto_dmInner_dmInner_tl_in_d_bits_size,
	auto_dmInner_dmInner_tl_in_d_bits_source,
	auto_dmInner_dmInner_tl_in_d_bits_data,
	auto_dmOuter_intsource_out_sync_0,
	io_debug_clock,
	io_debug_reset,
	io_ctrl_dmactive,
	io_ctrl_dmactiveAck,
	io_dmi_dmi_req_ready,
	io_dmi_dmi_req_valid,
	io_dmi_dmi_req_bits_addr,
	io_dmi_dmi_req_bits_data,
	io_dmi_dmi_req_bits_op,
	io_dmi_dmi_resp_ready,
	io_dmi_dmi_resp_valid,
	io_dmi_dmi_resp_bits_data,
	io_dmi_dmi_resp_bits_resp,
	io_dmi_dmiClock,
	io_dmi_dmiReset,
	io_hartIsInReset_0
);
	output wire auto_dmInner_dmInner_tl_in_a_ready;
	input auto_dmInner_dmInner_tl_in_a_valid;
	input [2:0] auto_dmInner_dmInner_tl_in_a_bits_opcode;
	input [2:0] auto_dmInner_dmInner_tl_in_a_bits_param;
	input [1:0] auto_dmInner_dmInner_tl_in_a_bits_size;
	input [7:0] auto_dmInner_dmInner_tl_in_a_bits_source;
	input [11:0] auto_dmInner_dmInner_tl_in_a_bits_address;
	input [3:0] auto_dmInner_dmInner_tl_in_a_bits_mask;
	input [31:0] auto_dmInner_dmInner_tl_in_a_bits_data;
	input auto_dmInner_dmInner_tl_in_a_bits_corrupt;
	input auto_dmInner_dmInner_tl_in_d_ready;
	output wire auto_dmInner_dmInner_tl_in_d_valid;
	output wire [2:0] auto_dmInner_dmInner_tl_in_d_bits_opcode;
	output wire [1:0] auto_dmInner_dmInner_tl_in_d_bits_size;
	output wire [7:0] auto_dmInner_dmInner_tl_in_d_bits_source;
	output wire [31:0] auto_dmInner_dmInner_tl_in_d_bits_data;
	output wire auto_dmOuter_intsource_out_sync_0;
	input io_debug_clock;
	input io_debug_reset;
	output wire io_ctrl_dmactive;
	input io_ctrl_dmactiveAck;
	output wire io_dmi_dmi_req_ready;
	input io_dmi_dmi_req_valid;
	input [6:0] io_dmi_dmi_req_bits_addr;
	input [31:0] io_dmi_dmi_req_bits_data;
	input [1:0] io_dmi_dmi_req_bits_op;
	input io_dmi_dmi_resp_ready;
	output wire io_dmi_dmi_resp_valid;
	output wire [31:0] io_dmi_dmi_resp_bits_data;
	output wire [1:0] io_dmi_dmi_resp_bits_resp;
	input io_dmi_dmiClock;
	input io_dmi_dmiReset;
	input io_hartIsInReset_0;
	wire [2:0] dmOuter_auto_asource_out_a_mem_0_opcode;
	wire [8:0] dmOuter_auto_asource_out_a_mem_0_address;
	wire [31:0] dmOuter_auto_asource_out_a_mem_0_data;
	wire dmOuter_auto_asource_out_a_ridx;
	wire dmOuter_auto_asource_out_a_widx;
	wire dmOuter_auto_asource_out_a_safe_ridx_valid;
	wire dmOuter_auto_asource_out_a_safe_widx_valid;
	wire dmOuter_auto_asource_out_a_safe_source_reset_n;
	wire dmOuter_auto_asource_out_a_safe_sink_reset_n;
	wire [2:0] dmOuter_auto_asource_out_d_mem_0_opcode;
	wire [1:0] dmOuter_auto_asource_out_d_mem_0_size;
	wire dmOuter_auto_asource_out_d_mem_0_source;
	wire [31:0] dmOuter_auto_asource_out_d_mem_0_data;
	wire dmOuter_auto_asource_out_d_ridx;
	wire dmOuter_auto_asource_out_d_widx;
	wire dmOuter_auto_asource_out_d_safe_ridx_valid;
	wire dmOuter_auto_asource_out_d_safe_widx_valid;
	wire dmOuter_auto_asource_out_d_safe_source_reset_n;
	wire dmOuter_auto_asource_out_d_safe_sink_reset_n;
	wire dmOuter_auto_intsource_out_sync_0;
	wire dmOuter_io_dmi_clock;
	wire dmOuter_io_dmi_reset;
	wire dmOuter_io_dmi_req_ready;
	wire dmOuter_io_dmi_req_valid;
	wire [6:0] dmOuter_io_dmi_req_bits_addr;
	wire [31:0] dmOuter_io_dmi_req_bits_data;
	wire [1:0] dmOuter_io_dmi_req_bits_op;
	wire dmOuter_io_dmi_resp_ready;
	wire dmOuter_io_dmi_resp_valid;
	wire [31:0] dmOuter_io_dmi_resp_bits_data;
	wire [1:0] dmOuter_io_dmi_resp_bits_resp;
	wire dmOuter_io_ctrl_dmactive;
	wire dmOuter_io_ctrl_dmactiveAck;
	wire dmOuter_io_innerCtrl_mem_0_resumereq;
	wire dmOuter_io_innerCtrl_mem_0_ackhavereset;
	wire dmOuter_io_innerCtrl_mem_0_hrmask_0;
	wire dmOuter_io_innerCtrl_ridx;
	wire dmOuter_io_innerCtrl_widx;
	wire dmOuter_io_innerCtrl_safe_ridx_valid;
	wire dmOuter_io_innerCtrl_safe_widx_valid;
	wire dmOuter_io_innerCtrl_safe_source_reset_n;
	wire dmOuter_io_innerCtrl_safe_sink_reset_n;
	wire dmOuter_io_hgDebugInt_0;
	wire [2:0] dmInner_auto_dmiXing_in_a_mem_0_opcode;
	wire [8:0] dmInner_auto_dmiXing_in_a_mem_0_address;
	wire [31:0] dmInner_auto_dmiXing_in_a_mem_0_data;
	wire dmInner_auto_dmiXing_in_a_ridx;
	wire dmInner_auto_dmiXing_in_a_widx;
	wire dmInner_auto_dmiXing_in_a_safe_ridx_valid;
	wire dmInner_auto_dmiXing_in_a_safe_widx_valid;
	wire dmInner_auto_dmiXing_in_a_safe_source_reset_n;
	wire dmInner_auto_dmiXing_in_a_safe_sink_reset_n;
	wire [2:0] dmInner_auto_dmiXing_in_d_mem_0_opcode;
	wire [1:0] dmInner_auto_dmiXing_in_d_mem_0_size;
	wire dmInner_auto_dmiXing_in_d_mem_0_source;
	wire [31:0] dmInner_auto_dmiXing_in_d_mem_0_data;
	wire dmInner_auto_dmiXing_in_d_ridx;
	wire dmInner_auto_dmiXing_in_d_widx;
	wire dmInner_auto_dmiXing_in_d_safe_ridx_valid;
	wire dmInner_auto_dmiXing_in_d_safe_widx_valid;
	wire dmInner_auto_dmiXing_in_d_safe_source_reset_n;
	wire dmInner_auto_dmiXing_in_d_safe_sink_reset_n;
	wire dmInner_auto_dmInner_tl_in_a_ready;
	wire dmInner_auto_dmInner_tl_in_a_valid;
	wire [2:0] dmInner_auto_dmInner_tl_in_a_bits_opcode;
	wire [2:0] dmInner_auto_dmInner_tl_in_a_bits_param;
	wire [1:0] dmInner_auto_dmInner_tl_in_a_bits_size;
	wire [7:0] dmInner_auto_dmInner_tl_in_a_bits_source;
	wire [11:0] dmInner_auto_dmInner_tl_in_a_bits_address;
	wire [3:0] dmInner_auto_dmInner_tl_in_a_bits_mask;
	wire [31:0] dmInner_auto_dmInner_tl_in_a_bits_data;
	wire dmInner_auto_dmInner_tl_in_a_bits_corrupt;
	wire dmInner_auto_dmInner_tl_in_d_ready;
	wire dmInner_auto_dmInner_tl_in_d_valid;
	wire [2:0] dmInner_auto_dmInner_tl_in_d_bits_opcode;
	wire [1:0] dmInner_auto_dmInner_tl_in_d_bits_size;
	wire [7:0] dmInner_auto_dmInner_tl_in_d_bits_source;
	wire [31:0] dmInner_auto_dmInner_tl_in_d_bits_data;
	wire dmInner_io_debug_clock;
	wire dmInner_io_debug_reset;
	wire dmInner_io_dmactive;
	wire dmInner_io_innerCtrl_mem_0_resumereq;
	wire dmInner_io_innerCtrl_mem_0_ackhavereset;
	wire dmInner_io_innerCtrl_mem_0_hrmask_0;
	wire dmInner_io_innerCtrl_ridx;
	wire dmInner_io_innerCtrl_widx;
	wire dmInner_io_innerCtrl_safe_ridx_valid;
	wire dmInner_io_innerCtrl_safe_widx_valid;
	wire dmInner_io_innerCtrl_safe_source_reset_n;
	wire dmInner_io_innerCtrl_safe_sink_reset_n;
	wire dmInner_io_hgDebugInt_0;
	wire dmInner_io_hartIsInReset_0;
	TLDebugModuleOuterAsync dmOuter(
		.auto_asource_out_a_mem_0_opcode(dmOuter_auto_asource_out_a_mem_0_opcode),
		.auto_asource_out_a_mem_0_address(dmOuter_auto_asource_out_a_mem_0_address),
		.auto_asource_out_a_mem_0_data(dmOuter_auto_asource_out_a_mem_0_data),
		.auto_asource_out_a_ridx(dmOuter_auto_asource_out_a_ridx),
		.auto_asource_out_a_widx(dmOuter_auto_asource_out_a_widx),
		.auto_asource_out_a_safe_ridx_valid(dmOuter_auto_asource_out_a_safe_ridx_valid),
		.auto_asource_out_a_safe_widx_valid(dmOuter_auto_asource_out_a_safe_widx_valid),
		.auto_asource_out_a_safe_source_reset_n(dmOuter_auto_asource_out_a_safe_source_reset_n),
		.auto_asource_out_a_safe_sink_reset_n(dmOuter_auto_asource_out_a_safe_sink_reset_n),
		.auto_asource_out_d_mem_0_opcode(dmOuter_auto_asource_out_d_mem_0_opcode),
		.auto_asource_out_d_mem_0_size(dmOuter_auto_asource_out_d_mem_0_size),
		.auto_asource_out_d_mem_0_source(dmOuter_auto_asource_out_d_mem_0_source),
		.auto_asource_out_d_mem_0_data(dmOuter_auto_asource_out_d_mem_0_data),
		.auto_asource_out_d_ridx(dmOuter_auto_asource_out_d_ridx),
		.auto_asource_out_d_widx(dmOuter_auto_asource_out_d_widx),
		.auto_asource_out_d_safe_ridx_valid(dmOuter_auto_asource_out_d_safe_ridx_valid),
		.auto_asource_out_d_safe_widx_valid(dmOuter_auto_asource_out_d_safe_widx_valid),
		.auto_asource_out_d_safe_source_reset_n(dmOuter_auto_asource_out_d_safe_source_reset_n),
		.auto_asource_out_d_safe_sink_reset_n(dmOuter_auto_asource_out_d_safe_sink_reset_n),
		.auto_intsource_out_sync_0(dmOuter_auto_intsource_out_sync_0),
		.io_dmi_clock(dmOuter_io_dmi_clock),
		.io_dmi_reset(dmOuter_io_dmi_reset),
		.io_dmi_req_ready(dmOuter_io_dmi_req_ready),
		.io_dmi_req_valid(dmOuter_io_dmi_req_valid),
		.io_dmi_req_bits_addr(dmOuter_io_dmi_req_bits_addr),
		.io_dmi_req_bits_data(dmOuter_io_dmi_req_bits_data),
		.io_dmi_req_bits_op(dmOuter_io_dmi_req_bits_op),
		.io_dmi_resp_ready(dmOuter_io_dmi_resp_ready),
		.io_dmi_resp_valid(dmOuter_io_dmi_resp_valid),
		.io_dmi_resp_bits_data(dmOuter_io_dmi_resp_bits_data),
		.io_dmi_resp_bits_resp(dmOuter_io_dmi_resp_bits_resp),
		.io_ctrl_dmactive(dmOuter_io_ctrl_dmactive),
		.io_ctrl_dmactiveAck(dmOuter_io_ctrl_dmactiveAck),
		.io_innerCtrl_mem_0_resumereq(dmOuter_io_innerCtrl_mem_0_resumereq),
		.io_innerCtrl_mem_0_ackhavereset(dmOuter_io_innerCtrl_mem_0_ackhavereset),
		.io_innerCtrl_mem_0_hrmask_0(dmOuter_io_innerCtrl_mem_0_hrmask_0),
		.io_innerCtrl_ridx(dmOuter_io_innerCtrl_ridx),
		.io_innerCtrl_widx(dmOuter_io_innerCtrl_widx),
		.io_innerCtrl_safe_ridx_valid(dmOuter_io_innerCtrl_safe_ridx_valid),
		.io_innerCtrl_safe_widx_valid(dmOuter_io_innerCtrl_safe_widx_valid),
		.io_innerCtrl_safe_source_reset_n(dmOuter_io_innerCtrl_safe_source_reset_n),
		.io_innerCtrl_safe_sink_reset_n(dmOuter_io_innerCtrl_safe_sink_reset_n),
		.io_hgDebugInt_0(dmOuter_io_hgDebugInt_0)
	);
	TLDebugModuleInnerAsync dmInner(
		.auto_dmiXing_in_a_mem_0_opcode(dmInner_auto_dmiXing_in_a_mem_0_opcode),
		.auto_dmiXing_in_a_mem_0_address(dmInner_auto_dmiXing_in_a_mem_0_address),
		.auto_dmiXing_in_a_mem_0_data(dmInner_auto_dmiXing_in_a_mem_0_data),
		.auto_dmiXing_in_a_ridx(dmInner_auto_dmiXing_in_a_ridx),
		.auto_dmiXing_in_a_widx(dmInner_auto_dmiXing_in_a_widx),
		.auto_dmiXing_in_a_safe_ridx_valid(dmInner_auto_dmiXing_in_a_safe_ridx_valid),
		.auto_dmiXing_in_a_safe_widx_valid(dmInner_auto_dmiXing_in_a_safe_widx_valid),
		.auto_dmiXing_in_a_safe_source_reset_n(dmInner_auto_dmiXing_in_a_safe_source_reset_n),
		.auto_dmiXing_in_a_safe_sink_reset_n(dmInner_auto_dmiXing_in_a_safe_sink_reset_n),
		.auto_dmiXing_in_d_mem_0_opcode(dmInner_auto_dmiXing_in_d_mem_0_opcode),
		.auto_dmiXing_in_d_mem_0_size(dmInner_auto_dmiXing_in_d_mem_0_size),
		.auto_dmiXing_in_d_mem_0_source(dmInner_auto_dmiXing_in_d_mem_0_source),
		.auto_dmiXing_in_d_mem_0_data(dmInner_auto_dmiXing_in_d_mem_0_data),
		.auto_dmiXing_in_d_ridx(dmInner_auto_dmiXing_in_d_ridx),
		.auto_dmiXing_in_d_widx(dmInner_auto_dmiXing_in_d_widx),
		.auto_dmiXing_in_d_safe_ridx_valid(dmInner_auto_dmiXing_in_d_safe_ridx_valid),
		.auto_dmiXing_in_d_safe_widx_valid(dmInner_auto_dmiXing_in_d_safe_widx_valid),
		.auto_dmiXing_in_d_safe_source_reset_n(dmInner_auto_dmiXing_in_d_safe_source_reset_n),
		.auto_dmiXing_in_d_safe_sink_reset_n(dmInner_auto_dmiXing_in_d_safe_sink_reset_n),
		.auto_dmInner_tl_in_a_ready(dmInner_auto_dmInner_tl_in_a_ready),
		.auto_dmInner_tl_in_a_valid(dmInner_auto_dmInner_tl_in_a_valid),
		.auto_dmInner_tl_in_a_bits_opcode(dmInner_auto_dmInner_tl_in_a_bits_opcode),
		.auto_dmInner_tl_in_a_bits_param(dmInner_auto_dmInner_tl_in_a_bits_param),
		.auto_dmInner_tl_in_a_bits_size(dmInner_auto_dmInner_tl_in_a_bits_size),
		.auto_dmInner_tl_in_a_bits_source(dmInner_auto_dmInner_tl_in_a_bits_source),
		.auto_dmInner_tl_in_a_bits_address(dmInner_auto_dmInner_tl_in_a_bits_address),
		.auto_dmInner_tl_in_a_bits_mask(dmInner_auto_dmInner_tl_in_a_bits_mask),
		.auto_dmInner_tl_in_a_bits_data(dmInner_auto_dmInner_tl_in_a_bits_data),
		.auto_dmInner_tl_in_a_bits_corrupt(dmInner_auto_dmInner_tl_in_a_bits_corrupt),
		.auto_dmInner_tl_in_d_ready(dmInner_auto_dmInner_tl_in_d_ready),
		.auto_dmInner_tl_in_d_valid(dmInner_auto_dmInner_tl_in_d_valid),
		.auto_dmInner_tl_in_d_bits_opcode(dmInner_auto_dmInner_tl_in_d_bits_opcode),
		.auto_dmInner_tl_in_d_bits_size(dmInner_auto_dmInner_tl_in_d_bits_size),
		.auto_dmInner_tl_in_d_bits_source(dmInner_auto_dmInner_tl_in_d_bits_source),
		.auto_dmInner_tl_in_d_bits_data(dmInner_auto_dmInner_tl_in_d_bits_data),
		.io_debug_clock(dmInner_io_debug_clock),
		.io_debug_reset(dmInner_io_debug_reset),
		.io_dmactive(dmInner_io_dmactive),
		.io_innerCtrl_mem_0_resumereq(dmInner_io_innerCtrl_mem_0_resumereq),
		.io_innerCtrl_mem_0_ackhavereset(dmInner_io_innerCtrl_mem_0_ackhavereset),
		.io_innerCtrl_mem_0_hrmask_0(dmInner_io_innerCtrl_mem_0_hrmask_0),
		.io_innerCtrl_ridx(dmInner_io_innerCtrl_ridx),
		.io_innerCtrl_widx(dmInner_io_innerCtrl_widx),
		.io_innerCtrl_safe_ridx_valid(dmInner_io_innerCtrl_safe_ridx_valid),
		.io_innerCtrl_safe_widx_valid(dmInner_io_innerCtrl_safe_widx_valid),
		.io_innerCtrl_safe_source_reset_n(dmInner_io_innerCtrl_safe_source_reset_n),
		.io_innerCtrl_safe_sink_reset_n(dmInner_io_innerCtrl_safe_sink_reset_n),
		.io_hgDebugInt_0(dmInner_io_hgDebugInt_0),
		.io_hartIsInReset_0(dmInner_io_hartIsInReset_0)
	);
	assign auto_dmInner_dmInner_tl_in_a_ready = dmInner_auto_dmInner_tl_in_a_ready;
	assign auto_dmInner_dmInner_tl_in_d_valid = dmInner_auto_dmInner_tl_in_d_valid;
	assign auto_dmInner_dmInner_tl_in_d_bits_opcode = dmInner_auto_dmInner_tl_in_d_bits_opcode;
	assign auto_dmInner_dmInner_tl_in_d_bits_size = dmInner_auto_dmInner_tl_in_d_bits_size;
	assign auto_dmInner_dmInner_tl_in_d_bits_source = dmInner_auto_dmInner_tl_in_d_bits_source;
	assign auto_dmInner_dmInner_tl_in_d_bits_data = dmInner_auto_dmInner_tl_in_d_bits_data;
	assign auto_dmOuter_intsource_out_sync_0 = dmOuter_auto_intsource_out_sync_0;
	assign io_ctrl_dmactive = dmOuter_io_ctrl_dmactive;
	assign io_dmi_dmi_req_ready = dmOuter_io_dmi_req_ready;
	assign io_dmi_dmi_resp_valid = dmOuter_io_dmi_resp_valid;
	assign io_dmi_dmi_resp_bits_data = dmOuter_io_dmi_resp_bits_data;
	assign io_dmi_dmi_resp_bits_resp = dmOuter_io_dmi_resp_bits_resp;
	assign dmOuter_auto_asource_out_a_ridx = dmInner_auto_dmiXing_in_a_ridx;
	assign dmOuter_auto_asource_out_a_safe_ridx_valid = dmInner_auto_dmiXing_in_a_safe_ridx_valid;
	assign dmOuter_auto_asource_out_a_safe_sink_reset_n = dmInner_auto_dmiXing_in_a_safe_sink_reset_n;
	assign dmOuter_auto_asource_out_d_mem_0_opcode = dmInner_auto_dmiXing_in_d_mem_0_opcode;
	assign dmOuter_auto_asource_out_d_mem_0_size = dmInner_auto_dmiXing_in_d_mem_0_size;
	assign dmOuter_auto_asource_out_d_mem_0_source = dmInner_auto_dmiXing_in_d_mem_0_source;
	assign dmOuter_auto_asource_out_d_mem_0_data = dmInner_auto_dmiXing_in_d_mem_0_data;
	assign dmOuter_auto_asource_out_d_widx = dmInner_auto_dmiXing_in_d_widx;
	assign dmOuter_auto_asource_out_d_safe_widx_valid = dmInner_auto_dmiXing_in_d_safe_widx_valid;
	assign dmOuter_auto_asource_out_d_safe_source_reset_n = dmInner_auto_dmiXing_in_d_safe_source_reset_n;
	assign dmOuter_io_dmi_clock = io_dmi_dmiClock;
	assign dmOuter_io_dmi_reset = io_dmi_dmiReset;
	assign dmOuter_io_dmi_req_valid = io_dmi_dmi_req_valid;
	assign dmOuter_io_dmi_req_bits_addr = io_dmi_dmi_req_bits_addr;
	assign dmOuter_io_dmi_req_bits_data = io_dmi_dmi_req_bits_data;
	assign dmOuter_io_dmi_req_bits_op = io_dmi_dmi_req_bits_op;
	assign dmOuter_io_dmi_resp_ready = io_dmi_dmi_resp_ready;
	assign dmOuter_io_ctrl_dmactiveAck = io_ctrl_dmactiveAck;
	assign dmOuter_io_innerCtrl_ridx = dmInner_io_innerCtrl_ridx;
	assign dmOuter_io_innerCtrl_safe_ridx_valid = dmInner_io_innerCtrl_safe_ridx_valid;
	assign dmOuter_io_innerCtrl_safe_sink_reset_n = dmInner_io_innerCtrl_safe_sink_reset_n;
	assign dmOuter_io_hgDebugInt_0 = dmInner_io_hgDebugInt_0;
	assign dmInner_auto_dmiXing_in_a_mem_0_opcode = dmOuter_auto_asource_out_a_mem_0_opcode;
	assign dmInner_auto_dmiXing_in_a_mem_0_address = dmOuter_auto_asource_out_a_mem_0_address;
	assign dmInner_auto_dmiXing_in_a_mem_0_data = dmOuter_auto_asource_out_a_mem_0_data;
	assign dmInner_auto_dmiXing_in_a_widx = dmOuter_auto_asource_out_a_widx;
	assign dmInner_auto_dmiXing_in_a_safe_widx_valid = dmOuter_auto_asource_out_a_safe_widx_valid;
	assign dmInner_auto_dmiXing_in_a_safe_source_reset_n = dmOuter_auto_asource_out_a_safe_source_reset_n;
	assign dmInner_auto_dmiXing_in_d_ridx = dmOuter_auto_asource_out_d_ridx;
	assign dmInner_auto_dmiXing_in_d_safe_ridx_valid = dmOuter_auto_asource_out_d_safe_ridx_valid;
	assign dmInner_auto_dmiXing_in_d_safe_sink_reset_n = dmOuter_auto_asource_out_d_safe_sink_reset_n;
	assign dmInner_auto_dmInner_tl_in_a_valid = auto_dmInner_dmInner_tl_in_a_valid;
	assign dmInner_auto_dmInner_tl_in_a_bits_opcode = auto_dmInner_dmInner_tl_in_a_bits_opcode;
	assign dmInner_auto_dmInner_tl_in_a_bits_param = auto_dmInner_dmInner_tl_in_a_bits_param;
	assign dmInner_auto_dmInner_tl_in_a_bits_size = auto_dmInner_dmInner_tl_in_a_bits_size;
	assign dmInner_auto_dmInner_tl_in_a_bits_source = auto_dmInner_dmInner_tl_in_a_bits_source;
	assign dmInner_auto_dmInner_tl_in_a_bits_address = auto_dmInner_dmInner_tl_in_a_bits_address;
	assign dmInner_auto_dmInner_tl_in_a_bits_mask = auto_dmInner_dmInner_tl_in_a_bits_mask;
	assign dmInner_auto_dmInner_tl_in_a_bits_data = auto_dmInner_dmInner_tl_in_a_bits_data;
	assign dmInner_auto_dmInner_tl_in_a_bits_corrupt = auto_dmInner_dmInner_tl_in_a_bits_corrupt;
	assign dmInner_auto_dmInner_tl_in_d_ready = auto_dmInner_dmInner_tl_in_d_ready;
	assign dmInner_io_debug_clock = io_debug_clock;
	assign dmInner_io_debug_reset = io_debug_reset;
	assign dmInner_io_dmactive = dmOuter_io_ctrl_dmactive;
	assign dmInner_io_innerCtrl_mem_0_resumereq = dmOuter_io_innerCtrl_mem_0_resumereq;
	assign dmInner_io_innerCtrl_mem_0_ackhavereset = dmOuter_io_innerCtrl_mem_0_ackhavereset;
	assign dmInner_io_innerCtrl_mem_0_hrmask_0 = dmOuter_io_innerCtrl_mem_0_hrmask_0;
	assign dmInner_io_innerCtrl_widx = dmOuter_io_innerCtrl_widx;
	assign dmInner_io_innerCtrl_safe_widx_valid = dmOuter_io_innerCtrl_safe_widx_valid;
	assign dmInner_io_innerCtrl_safe_source_reset_n = dmOuter_io_innerCtrl_safe_source_reset_n;
	assign dmInner_io_hartIsInReset_0 = io_hartIsInReset_0;
endmodule
module BundleBridgeNexus_13 (auto_out);
	output wire auto_out;
	wire outputs_0 = 1'h0;
	assign auto_out = outputs_0;
endmodule
module AsyncResetRegVec_w2_i0 (
	clock,
	reset,
	io_d,
	io_q
);
	input clock;
	input reset;
	input [1:0] io_d;
	output wire [1:0] io_q;
	reg [1:0] reg_;
	assign io_q = reg_;
	always @(posedge clock or posedge reset)
		if (reset)
			reg_ <= 2'h0;
		else
			reg_ <= io_d;
endmodule
module IntSyncCrossingSource_5 (
	clock,
	reset,
	auto_in_0,
	auto_in_1,
	auto_out_sync_0,
	auto_out_sync_1
);
	input clock;
	input reset;
	input auto_in_0;
	input auto_in_1;
	output wire auto_out_sync_0;
	output wire auto_out_sync_1;
	wire reg__clock;
	wire reg__reset;
	wire [1:0] reg__io_d;
	wire [1:0] reg__io_q;
	AsyncResetRegVec_w2_i0 reg_(
		.clock(reg__clock),
		.reset(reg__reset),
		.io_d(reg__io_d),
		.io_q(reg__io_q)
	);
	assign auto_out_sync_0 = reg__io_q[0];
	assign auto_out_sync_1 = reg__io_q[1];
	assign reg__clock = clock;
	assign reg__reset = reset;
	assign reg__io_d = {auto_in_1, auto_in_0};
endmodule
module TLMonitor_43 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [1:0] io_in_a_bits_size;
	input [7:0] io_in_a_bits_source;
	input [16:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [1:0] io_in_d_bits_size;
	input [7:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_4 = io_in_a_bits_source <= 8'h9f;
	wire [4:0] _is_aligned_mask_T_1 = 5'h03 << io_in_a_bits_size;
	wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0];
	wire [16:0] _GEN_71 = {15'd0, is_aligned_mask};
	wire [16:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 17'h00000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 2'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_10 = ~_source_ok_T_4;
	wire _T_20 = io_in_a_bits_opcode == 3'h6;
	wire [16:0] _T_33 = io_in_a_bits_address ^ 17'h10000;
	wire [17:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [17:0] _T_36 = $signed(_T_34) & -18'sh10000;
	wire _T_37 = $signed(_T_36) == 18'sh00000;
	wire _T_69 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_73 = ~io_in_a_bits_mask;
	wire _T_74 = _T_73 == 4'h0;
	wire _T_78 = ~io_in_a_bits_corrupt;
	wire _T_82 = io_in_a_bits_opcode == 3'h7;
	wire _T_135 = io_in_a_bits_param != 3'h0;
	wire _T_148 = io_in_a_bits_opcode == 3'h4;
	wire _T_164 = io_in_a_bits_size <= 2'h2;
	wire _T_172 = _T_164 & _T_37;
	wire _T_183 = io_in_a_bits_param == 3'h0;
	wire _T_187 = io_in_a_bits_mask == mask;
	wire _T_195 = io_in_a_bits_opcode == 3'h0;
	wire _T_233 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_267 = ~mask;
	wire [3:0] _T_268 = io_in_a_bits_mask & _T_267;
	wire _T_269 = _T_268 == 4'h0;
	wire _T_273 = io_in_a_bits_opcode == 3'h2;
	wire _T_303 = io_in_a_bits_param <= 3'h4;
	wire _T_311 = io_in_a_bits_opcode == 3'h3;
	wire _T_341 = io_in_a_bits_param <= 3'h3;
	wire _T_349 = io_in_a_bits_opcode == 3'h5;
	wire _T_379 = io_in_a_bits_param <= 3'h1;
	wire _source_ok_T_10 = io_in_d_bits_source <= 8'h9f;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [1:0] size;
	reg [7:0] source;
	reg [16:0] address;
	wire _T_537 = io_in_a_valid & ~a_first;
	wire _T_538 = io_in_a_bits_opcode == opcode;
	wire _T_542 = io_in_a_bits_param == param;
	wire _T_546 = io_in_a_bits_size == size;
	wire _T_550 = io_in_a_bits_source == source;
	wire _T_554 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [1:0] size_1;
	reg [7:0] source_1;
	wire _T_561 = io_in_d_valid & ~d_first;
	wire _T_570 = io_in_d_bits_size == size_1;
	wire _T_574 = io_in_d_bits_source == source_1;
	reg [159:0] inflight;
	reg [639:0] inflight_opcodes;
	reg [639:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [10:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [639:0] _GEN_73 = {624'd0, _a_opcode_lookup_T_5};
	wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [639:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[639:1]};
	wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [639:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[639:1]};
	wire _T_588 = io_in_a_valid & a_first_1;
	wire [255:0] _a_set_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_a_bits_source;
	wire _T_591 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1;
	wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [10:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [2050:0] _GEN_1 = {2047'd0, a_opcodes_set_interm};
	wire [2050:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? _a_sizes_set_interm_T_1 : 3'h0);
	wire [2049:0] _GEN_2 = {2047'd0, a_sizes_set_interm};
	wire [2049:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [159:0] _T_593 = inflight >> io_in_a_bits_source;
	wire _T_595 = ~_T_593[0];
	wire [255:0] _GEN_16 = (a_first_done & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2050:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 2051'h0);
	wire [2049:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 2050'h0);
	wire _T_599 = io_in_d_valid & d_first_1;
	wire [255:0] _d_clr_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_d_bits_source;
	wire [2062:0] _GEN_3 = {2047'd0, _a_opcode_lookup_T_5};
	wire [2062:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [255:0] _GEN_22 = (d_first_done & d_first_1 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_23 = (d_first_done & d_first_1 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_588 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [159:0] _T_612 = inflight >> io_in_d_bits_source;
	wire _T_614 = _T_612[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_619 = 3'h1 == _GEN_40;
	wire _T_620 = (3'h1 == _GEN_32) | _T_619;
	wire _T_624 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_631 = 3'h1 == _GEN_56;
	wire _T_632 = (3'h1 == _GEN_48) | _T_631;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {2'd0, io_in_d_bits_size};
	wire _T_636 = _GEN_82 == a_size_lookup;
	wire _T_644 = ((_T_599 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2;
	wire _T_648 = ~io_in_d_ready | io_in_a_ready;
	wire [159:0] a_set = _GEN_16[159:0];
	wire [159:0] _inflight_T = inflight | a_set;
	wire [159:0] d_clr = _GEN_22[159:0];
	wire [159:0] _inflight_T_1 = ~d_clr;
	wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [639:0] a_opcodes_set = _GEN_19[639:0];
	wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [639:0] d_opcodes_clr = _GEN_23[639:0];
	wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [639:0] a_sizes_set = _GEN_20[639:0];
	wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_657 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			param <= io_in_a_bits_param;
		if (a_first_done & a_first)
			size <= io_in_a_bits_size;
		if (a_first_done & a_first)
			source <= io_in_a_bits_source;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 160'h0000000000000000000000000000000000000000;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 640'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 640'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
	end
endmodule
module TLROM (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [1:0] auto_in_a_bits_size;
	input [7:0] auto_in_a_bits_source;
	input [16:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [1:0] auto_in_d_bits_size;
	output wire [7:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [1:0] monitor_io_in_a_bits_size;
	wire [7:0] monitor_io_in_a_bits_source;
	wire [16:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [1:0] monitor_io_in_d_bits_size;
	wire [7:0] monitor_io_in_d_bits_source;
	wire [9:0] index = auto_in_a_bits_address[11:2];
	wire [3:0] high = auto_in_a_bits_address[15:12];
	wire [31:0] _GEN_1 = (10'h001 == index ? 32'hf1402573 : 32'h020005b7);
	wire [31:0] _GEN_2 = (10'h002 == index ? 32'h00050463 : _GEN_1);
	wire [31:0] _GEN_3 = (10'h003 == index ? 32'h0780006f : _GEN_2);
	wire [31:0] _GEN_4 = (10'h004 == index ? 32'h00458613 : _GEN_3);
	wire [31:0] _GEN_5 = (10'h005 == index ? 32'h00100693 : _GEN_4);
	wire [31:0] _GEN_6 = (10'h006 == index ? 32'h00d62023 : _GEN_5);
	wire [31:0] _GEN_7 = (10'h007 == index ? 32'h00460613 : _GEN_6);
	wire [31:0] _GEN_8 = (10'h008 == index ? 32'hffc62683 : _GEN_7);
	wire [31:0] _GEN_9 = (10'h009 == index ? 32'hfe069ae3 : _GEN_8);
	wire [31:0] _GEN_10 = (10'h00a == index ? 32'h06c0006f : _GEN_9);
	wire [31:0] _GEN_11 = (10'h00b == index ? 32'h00000000 : _GEN_10);
	wire [31:0] _GEN_12 = (10'h00c == index ? 32'h00000000 : _GEN_11);
	wire [31:0] _GEN_13 = (10'h00d == index ? 32'h00000000 : _GEN_12);
	wire [31:0] _GEN_14 = (10'h00e == index ? 32'h00000000 : _GEN_13);
	wire [31:0] _GEN_15 = (10'h00f == index ? 32'h00000000 : _GEN_14);
	wire [31:0] _GEN_16 = (10'h010 == index ? 32'h00000517 : _GEN_15);
	wire [31:0] _GEN_17 = (10'h011 == index ? 32'hfc050513 : _GEN_16);
	wire [31:0] _GEN_18 = (10'h012 == index ? 32'h30551073 : _GEN_17);
	wire [31:0] _GEN_19 = (10'h013 == index ? 32'h301022f3 : _GEN_18);
	wire [31:0] _GEN_20 = (10'h014 == index ? 32'h4122d293 : _GEN_19);
	wire [31:0] _GEN_21 = (10'h015 == index ? 32'h0012f293 : _GEN_20);
	wire [31:0] _GEN_22 = (10'h016 == index ? 32'h00028463 : _GEN_21);
	wire [31:0] _GEN_23 = (10'h017 == index ? 32'h30301073 : _GEN_22);
	wire [31:0] _GEN_24 = (10'h018 == index ? 32'h00800513 : _GEN_23);
	wire [31:0] _GEN_25 = (10'h019 == index ? 32'h30451073 : _GEN_24);
	wire [31:0] _GEN_26 = (10'h01a == index ? 32'h30052073 : _GEN_25);
	wire [31:0] _GEN_27 = (10'h01b == index ? 32'h10500073 : _GEN_26);
	wire [31:0] _GEN_28 = (10'h01c == index ? 32'hffdff06f : _GEN_27);
	wire [31:0] _GEN_29 = (10'h01d == index ? 32'h00000000 : _GEN_28);
	wire [31:0] _GEN_30 = (10'h01e == index ? 32'h00000000 : _GEN_29);
	wire [31:0] _GEN_31 = (10'h01f == index ? 32'h00000000 : _GEN_30);
	wire [31:0] _GEN_32 = (10'h020 == index ? 32'hfc1ff06f : _GEN_31);
	wire [31:0] _GEN_33 = (10'h021 == index ? 32'h0005a283 : _GEN_32);
	wire [31:0] _GEN_34 = (10'h022 == index ? 32'hfe029ee3 : _GEN_33);
	wire [31:0] _GEN_35 = (10'h023 == index ? 32'h00251513 : _GEN_34);
	wire [31:0] _GEN_36 = (10'h024 == index ? 32'h00b505b3 : _GEN_35);
	wire [31:0] _GEN_37 = (10'h025 == index ? 32'h0005a023 : _GEN_36);
	wire [31:0] _GEN_38 = (10'h026 == index ? 32'h00004537 : _GEN_37);
	wire [31:0] _GEN_39 = (10'h027 == index ? 32'h00052503 : _GEN_38);
	wire [31:0] _GEN_40 = (10'h028 == index ? 32'h34151073 : _GEN_39);
	wire [31:0] _GEN_41 = (10'h029 == index ? 32'hf1402573 : _GEN_40);
	wire [31:0] _GEN_42 = (10'h02a == index ? 32'h00000597 : _GEN_41);
	wire [31:0] _GEN_43 = (10'h02b == index ? 32'h01858593 : _GEN_42);
	wire [31:0] _GEN_44 = (10'h02c == index ? 32'h08000613 : _GEN_43);
	wire [31:0] _GEN_45 = (10'h02d == index ? 32'h30063073 : _GEN_44);
	wire [31:0] _GEN_46 = (10'h02e == index ? 32'h30200073 : _GEN_45);
	wire [31:0] _GEN_47 = (10'h02f == index ? 32'h00000013 : _GEN_46);
	wire [31:0] _GEN_48 = (10'h030 == index ? 32'hedfe0dd0 : _GEN_47);
	wire [31:0] _GEN_49 = (10'h031 == index ? 32'h2b0a0000 : _GEN_48);
	wire [31:0] _GEN_50 = (10'h032 == index ? 32'h38000000 : _GEN_49);
	wire [31:0] _GEN_51 = (10'h033 == index ? 32'h74080000 : _GEN_50);
	wire [31:0] _GEN_52 = (10'h034 == index ? 32'h28000000 : _GEN_51);
	wire [31:0] _GEN_53 = (10'h035 == index ? 32'h11000000 : _GEN_52);
	wire [31:0] _GEN_54 = (10'h036 == index ? 32'h10000000 : _GEN_53);
	wire [31:0] _GEN_55 = (10'h037 == index ? 32'h00000000 : _GEN_54);
	wire [31:0] _GEN_56 = (10'h038 == index ? 32'hb7010000 : _GEN_55);
	wire [31:0] _GEN_57 = (10'h039 == index ? 32'h3c080000 : _GEN_56);
	wire [31:0] _GEN_58 = (10'h03a == index ? 32'h00000000 : _GEN_57);
	wire [31:0] _GEN_59 = (10'h03b == index ? 32'h00000000 : _GEN_58);
	wire [31:0] _GEN_60 = (10'h03c == index ? 32'h00000000 : _GEN_59);
	wire [31:0] _GEN_61 = (10'h03d == index ? 32'h00000000 : _GEN_60);
	wire [31:0] _GEN_62 = (10'h03e == index ? 32'h01000000 : _GEN_61);
	wire [31:0] _GEN_63 = (10'h03f == index ? 32'h00000000 : _GEN_62);
	wire [31:0] _GEN_64 = (10'h040 == index ? 32'h03000000 : _GEN_63);
	wire [31:0] _GEN_65 = (10'h041 == index ? 32'h04000000 : _GEN_64);
	wire [31:0] _GEN_66 = (10'h042 == index ? 32'h00000000 : _GEN_65);
	wire [31:0] _GEN_67 = (10'h043 == index ? 32'h01000000 : _GEN_66);
	wire [31:0] _GEN_68 = (10'h044 == index ? 32'h03000000 : _GEN_67);
	wire [31:0] _GEN_69 = (10'h045 == index ? 32'h04000000 : _GEN_68);
	wire [31:0] _GEN_70 = (10'h046 == index ? 32'h0f000000 : _GEN_69);
	wire [31:0] _GEN_71 = (10'h047 == index ? 32'h01000000 : _GEN_70);
	wire [31:0] _GEN_72 = (10'h048 == index ? 32'h03000000 : _GEN_71);
	wire [31:0] _GEN_73 = (10'h049 == index ? 32'h21000000 : _GEN_72);
	wire [31:0] _GEN_74 = (10'h04a == index ? 32'h1b000000 : _GEN_73);
	wire [31:0] _GEN_75 = (10'h04b == index ? 32'h65657266 : _GEN_74);
	wire [31:0] _GEN_76 = (10'h04c == index ? 32'h70696863 : _GEN_75);
	wire [31:0] _GEN_77 = (10'h04d == index ? 32'h6f722c73 : _GEN_76);
	wire [31:0] _GEN_78 = (10'h04e == index ? 32'h74656b63 : _GEN_77);
	wire [31:0] _GEN_79 = (10'h04f == index ? 32'h70696863 : _GEN_78);
	wire [31:0] _GEN_80 = (10'h050 == index ? 32'h6b6e752d : _GEN_79);
	wire [31:0] _GEN_81 = (10'h051 == index ? 32'h6e776f6e : _GEN_80);
	wire [31:0] _GEN_82 = (10'h052 == index ? 32'h7665642d : _GEN_81);
	wire [31:0] _GEN_83 = (10'h053 == index ? 32'h00000000 : _GEN_82);
	wire [31:0] _GEN_84 = (10'h054 == index ? 32'h03000000 : _GEN_83);
	wire [31:0] _GEN_85 = (10'h055 == index ? 32'h1d000000 : _GEN_84);
	wire [31:0] _GEN_86 = (10'h056 == index ? 32'h26000000 : _GEN_85);
	wire [31:0] _GEN_87 = (10'h057 == index ? 32'h65657266 : _GEN_86);
	wire [31:0] _GEN_88 = (10'h058 == index ? 32'h70696863 : _GEN_87);
	wire [31:0] _GEN_89 = (10'h059 == index ? 32'h6f722c73 : _GEN_88);
	wire [31:0] _GEN_90 = (10'h05a == index ? 32'h74656b63 : _GEN_89);
	wire [31:0] _GEN_91 = (10'h05b == index ? 32'h70696863 : _GEN_90);
	wire [31:0] _GEN_92 = (10'h05c == index ? 32'h6b6e752d : _GEN_91);
	wire [31:0] _GEN_93 = (10'h05d == index ? 32'h6e776f6e : _GEN_92);
	wire [31:0] _GEN_94 = (10'h05e == index ? 32'h00000000 : _GEN_93);
	wire [31:0] _GEN_95 = (10'h05f == index ? 32'h01000000 : _GEN_94);
	wire [31:0] _GEN_96 = (10'h060 == index ? 32'h61696c61 : _GEN_95);
	wire [31:0] _GEN_97 = (10'h061 == index ? 32'h00736573 : _GEN_96);
	wire [31:0] _GEN_98 = (10'h062 == index ? 32'h03000000 : _GEN_97);
	wire [31:0] _GEN_99 = (10'h063 == index ? 32'h15000000 : _GEN_98);
	wire [31:0] _GEN_100 = (10'h064 == index ? 32'h2c000000 : _GEN_99);
	wire [31:0] _GEN_101 = (10'h065 == index ? 32'h636f732f : _GEN_100);
	wire [31:0] _GEN_102 = (10'h066 == index ? 32'h7265732f : _GEN_101);
	wire [31:0] _GEN_103 = (10'h067 == index ? 32'h406c6169 : _GEN_102);
	wire [31:0] _GEN_104 = (10'h068 == index ? 32'h30303435 : _GEN_103);
	wire [31:0] _GEN_105 = (10'h069 == index ? 32'h30303030 : _GEN_104);
	wire [31:0] _GEN_106 = (10'h06a == index ? 32'h00000000 : _GEN_105);
	wire [31:0] _GEN_107 = (10'h06b == index ? 32'h02000000 : _GEN_106);
	wire [31:0] _GEN_108 = (10'h06c == index ? 32'h01000000 : _GEN_107);
	wire [31:0] _GEN_109 = (10'h06d == index ? 32'h73757063 : _GEN_108);
	wire [31:0] _GEN_110 = (10'h06e == index ? 32'h00000000 : _GEN_109);
	wire [31:0] _GEN_111 = (10'h06f == index ? 32'h03000000 : _GEN_110);
	wire [31:0] _GEN_112 = (10'h070 == index ? 32'h04000000 : _GEN_111);
	wire [31:0] _GEN_113 = (10'h071 == index ? 32'h00000000 : _GEN_112);
	wire [31:0] _GEN_114 = (10'h072 == index ? 32'h01000000 : _GEN_113);
	wire [31:0] _GEN_115 = (10'h073 == index ? 32'h03000000 : _GEN_114);
	wire [31:0] _GEN_116 = (10'h074 == index ? 32'h04000000 : _GEN_115);
	wire [31:0] _GEN_117 = (10'h075 == index ? 32'h0f000000 : _GEN_116);
	wire [31:0] _GEN_118 = (10'h076 == index ? 32'h00000000 : _GEN_117);
	wire [31:0] _GEN_119 = (10'h077 == index ? 32'h03000000 : _GEN_118);
	wire [31:0] _GEN_120 = (10'h078 == index ? 32'h04000000 : _GEN_119);
	wire [31:0] _GEN_121 = (10'h079 == index ? 32'h34000000 : _GEN_120);
	wire [31:0] _GEN_122 = (10'h07a == index ? 32'h40420f00 : _GEN_121);
	wire [31:0] _GEN_123 = (10'h07b == index ? 32'h01000000 : _GEN_122);
	wire [31:0] _GEN_124 = (10'h07c == index ? 32'h40757063 : _GEN_123);
	wire [31:0] _GEN_125 = (10'h07d == index ? 32'h00000030 : _GEN_124);
	wire [31:0] _GEN_126 = (10'h07e == index ? 32'h03000000 : _GEN_125);
	wire [31:0] _GEN_127 = (10'h07f == index ? 32'h04000000 : _GEN_126);
	wire [31:0] _GEN_128 = (10'h080 == index ? 32'h47000000 : _GEN_127);
	wire [31:0] _GEN_129 = (10'h081 == index ? 32'h00000000 : _GEN_128);
	wire [31:0] _GEN_130 = (10'h082 == index ? 32'h03000000 : _GEN_129);
	wire [31:0] _GEN_131 = (10'h083 == index ? 32'h15000000 : _GEN_130);
	wire [31:0] _GEN_132 = (10'h084 == index ? 32'h1b000000 : _GEN_131);
	wire [31:0] _GEN_133 = (10'h085 == index ? 32'h69666973 : _GEN_132);
	wire [31:0] _GEN_134 = (10'h086 == index ? 32'h722c6576 : _GEN_133);
	wire [31:0] _GEN_135 = (10'h087 == index ? 32'h656b636f : _GEN_134);
	wire [31:0] _GEN_136 = (10'h088 == index ? 32'h72003074 : _GEN_135);
	wire [31:0] _GEN_137 = (10'h089 == index ? 32'h76637369 : _GEN_136);
	wire [31:0] _GEN_138 = (10'h08a == index ? 32'h00000000 : _GEN_137);
	wire [31:0] _GEN_139 = (10'h08b == index ? 32'h03000000 : _GEN_138);
	wire [31:0] _GEN_140 = (10'h08c == index ? 32'h04000000 : _GEN_139);
	wire [31:0] _GEN_141 = (10'h08d == index ? 32'h57000000 : _GEN_140);
	wire [31:0] _GEN_142 = (10'h08e == index ? 32'h00757063 : _GEN_141);
	wire [31:0] _GEN_143 = (10'h08f == index ? 32'h03000000 : _GEN_142);
	wire [31:0] _GEN_144 = (10'h090 == index ? 32'h04000000 : _GEN_143);
	wire [31:0] _GEN_145 = (10'h091 == index ? 32'h63000000 : _GEN_144);
	wire [31:0] _GEN_146 = (10'h092 == index ? 32'h01000000 : _GEN_145);
	wire [31:0] _GEN_147 = (10'h093 == index ? 32'h03000000 : _GEN_146);
	wire [31:0] _GEN_148 = (10'h094 == index ? 32'h04000000 : _GEN_147);
	wire [31:0] _GEN_149 = (10'h095 == index ? 32'h82000000 : _GEN_148);
	wire [31:0] _GEN_150 = (10'h096 == index ? 32'h40000000 : _GEN_149);
	wire [31:0] _GEN_151 = (10'h097 == index ? 32'h03000000 : _GEN_150);
	wire [31:0] _GEN_152 = (10'h098 == index ? 32'h04000000 : _GEN_151);
	wire [31:0] _GEN_153 = (10'h099 == index ? 32'h95000000 : _GEN_152);
	wire [31:0] _GEN_154 = (10'h09a == index ? 32'h40000000 : _GEN_153);
	wire [31:0] _GEN_155 = (10'h09b == index ? 32'h03000000 : _GEN_154);
	wire [31:0] _GEN_156 = (10'h09c == index ? 32'h04000000 : _GEN_155);
	wire [31:0] _GEN_157 = (10'h09d == index ? 32'ha2000000 : _GEN_156);
	wire [31:0] _GEN_158 = (10'h09e == index ? 32'h00100000 : _GEN_157);
	wire [31:0] _GEN_159 = (10'h09f == index ? 32'h03000000 : _GEN_158);
	wire [31:0] _GEN_160 = (10'h0a0 == index ? 32'h04000000 : _GEN_159);
	wire [31:0] _GEN_161 = (10'h0a1 == index ? 32'haf000000 : _GEN_160);
	wire [31:0] _GEN_162 = (10'h0a2 == index ? 32'h00000000 : _GEN_161);
	wire [31:0] _GEN_163 = (10'h0a3 == index ? 32'h03000000 : _GEN_162);
	wire [31:0] _GEN_164 = (10'h0a4 == index ? 32'h09000000 : _GEN_163);
	wire [31:0] _GEN_165 = (10'h0a5 == index ? 32'hb3000000 : _GEN_164);
	wire [31:0] _GEN_166 = (10'h0a6 == index ? 32'h32337672 : _GEN_165);
	wire [31:0] _GEN_167 = (10'h0a7 == index ? 32'h63616d69 : _GEN_166);
	wire [31:0] _GEN_168 = (10'h0a8 == index ? 32'h00000000 : _GEN_167);
	wire [31:0] _GEN_169 = (10'h0a9 == index ? 32'h03000000 : _GEN_168);
	wire [31:0] _GEN_170 = (10'h0aa == index ? 32'h04000000 : _GEN_169);
	wire [31:0] _GEN_171 = (10'h0ab == index ? 32'hbd000000 : _GEN_170);
	wire [31:0] _GEN_172 = (10'h0ac == index ? 32'h04000000 : _GEN_171);
	wire [31:0] _GEN_173 = (10'h0ad == index ? 32'h03000000 : _GEN_172);
	wire [31:0] _GEN_174 = (10'h0ae == index ? 32'h04000000 : _GEN_173);
	wire [31:0] _GEN_175 = (10'h0af == index ? 32'hd2000000 : _GEN_174);
	wire [31:0] _GEN_176 = (10'h0b0 == index ? 32'h08000000 : _GEN_175);
	wire [31:0] _GEN_177 = (10'h0b1 == index ? 32'h03000000 : _GEN_176);
	wire [31:0] _GEN_178 = (10'h0b2 == index ? 32'h04000000 : _GEN_177);
	wire [31:0] _GEN_179 = (10'h0b3 == index ? 32'he3000000 : _GEN_178);
	wire [31:0] _GEN_180 = (10'h0b4 == index ? 32'h01000000 : _GEN_179);
	wire [31:0] _GEN_181 = (10'h0b5 == index ? 32'h03000000 : _GEN_180);
	wire [31:0] _GEN_182 = (10'h0b6 == index ? 32'h05000000 : _GEN_181);
	wire [31:0] _GEN_183 = (10'h0b7 == index ? 32'hef000000 : _GEN_182);
	wire [31:0] _GEN_184 = (10'h0b8 == index ? 32'h79616b6f : _GEN_183);
	wire [31:0] _GEN_185 = (10'h0b9 == index ? 32'h00000000 : _GEN_184);
	wire [31:0] _GEN_186 = (10'h0ba == index ? 32'h03000000 : _GEN_185);
	wire [31:0] _GEN_187 = (10'h0bb == index ? 32'h04000000 : _GEN_186);
	wire [31:0] _GEN_188 = (10'h0bc == index ? 32'h34000000 : _GEN_187);
	wire [31:0] _GEN_189 = (10'h0bd == index ? 32'h40420f00 : _GEN_188);
	wire [31:0] _GEN_190 = (10'h0be == index ? 32'h01000000 : _GEN_189);
	wire [31:0] _GEN_191 = (10'h0bf == index ? 32'h65746e69 : _GEN_190);
	wire [31:0] _GEN_192 = (10'h0c0 == index ? 32'h70757272 : _GEN_191);
	wire [31:0] _GEN_193 = (10'h0c1 == index ? 32'h6f632d74 : _GEN_192);
	wire [31:0] _GEN_194 = (10'h0c2 == index ? 32'h6f72746e : _GEN_193);
	wire [31:0] _GEN_195 = (10'h0c3 == index ? 32'h72656c6c : _GEN_194);
	wire [31:0] _GEN_196 = (10'h0c4 == index ? 32'h00000000 : _GEN_195);
	wire [31:0] _GEN_197 = (10'h0c5 == index ? 32'h03000000 : _GEN_196);
	wire [31:0] _GEN_198 = (10'h0c6 == index ? 32'h04000000 : _GEN_197);
	wire [31:0] _GEN_199 = (10'h0c7 == index ? 32'hf6000000 : _GEN_198);
	wire [31:0] _GEN_200 = (10'h0c8 == index ? 32'h01000000 : _GEN_199);
	wire [31:0] _GEN_201 = (10'h0c9 == index ? 32'h03000000 : _GEN_200);
	wire [31:0] _GEN_202 = (10'h0ca == index ? 32'h0f000000 : _GEN_201);
	wire [31:0] _GEN_203 = (10'h0cb == index ? 32'h1b000000 : _GEN_202);
	wire [31:0] _GEN_204 = (10'h0cc == index ? 32'h63736972 : _GEN_203);
	wire [31:0] _GEN_205 = (10'h0cd == index ? 32'h70632c76 : _GEN_204);
	wire [31:0] _GEN_206 = (10'h0ce == index ? 32'h6e692d75 : _GEN_205);
	wire [31:0] _GEN_207 = (10'h0cf == index ? 32'h00006374 : _GEN_206);
	wire [31:0] _GEN_208 = (10'h0d0 == index ? 32'h03000000 : _GEN_207);
	wire [31:0] _GEN_209 = (10'h0d1 == index ? 32'h00000000 : _GEN_208);
	wire [31:0] _GEN_210 = (10'h0d2 == index ? 32'h07010000 : _GEN_209);
	wire [31:0] _GEN_211 = (10'h0d3 == index ? 32'h03000000 : _GEN_210);
	wire [31:0] _GEN_212 = (10'h0d4 == index ? 32'h04000000 : _GEN_211);
	wire [31:0] _GEN_213 = (10'h0d5 == index ? 32'h1c010000 : _GEN_212);
	wire [31:0] _GEN_214 = (10'h0d6 == index ? 32'h02000000 : _GEN_213);
	wire [31:0] _GEN_215 = (10'h0d7 == index ? 32'h02000000 : _GEN_214);
	wire [31:0] _GEN_216 = (10'h0d8 == index ? 32'h02000000 : _GEN_215);
	wire [31:0] _GEN_217 = (10'h0d9 == index ? 32'h02000000 : _GEN_216);
	wire [31:0] _GEN_218 = (10'h0da == index ? 32'h01000000 : _GEN_217);
	wire [31:0] _GEN_219 = (10'h0db == index ? 32'h66697468 : _GEN_218);
	wire [31:0] _GEN_220 = (10'h0dc == index ? 32'h00000000 : _GEN_219);
	wire [31:0] _GEN_221 = (10'h0dd == index ? 32'h03000000 : _GEN_220);
	wire [31:0] _GEN_222 = (10'h0de == index ? 32'h0a000000 : _GEN_221);
	wire [31:0] _GEN_223 = (10'h0df == index ? 32'h1b000000 : _GEN_222);
	wire [31:0] _GEN_224 = (10'h0e0 == index ? 32'h2c626375 : _GEN_223);
	wire [31:0] _GEN_225 = (10'h0e1 == index ? 32'h66697468 : _GEN_224);
	wire [31:0] _GEN_226 = (10'h0e2 == index ? 32'h00000030 : _GEN_225);
	wire [31:0] _GEN_227 = (10'h0e3 == index ? 32'h02000000 : _GEN_226);
	wire [31:0] _GEN_228 = (10'h0e4 == index ? 32'h01000000 : _GEN_227);
	wire [31:0] _GEN_229 = (10'h0e5 == index ? 32'h00636f73 : _GEN_228);
	wire [31:0] _GEN_230 = (10'h0e6 == index ? 32'h03000000 : _GEN_229);
	wire [31:0] _GEN_231 = (10'h0e7 == index ? 32'h04000000 : _GEN_230);
	wire [31:0] _GEN_232 = (10'h0e8 == index ? 32'h00000000 : _GEN_231);
	wire [31:0] _GEN_233 = (10'h0e9 == index ? 32'h01000000 : _GEN_232);
	wire [31:0] _GEN_234 = (10'h0ea == index ? 32'h03000000 : _GEN_233);
	wire [31:0] _GEN_235 = (10'h0eb == index ? 32'h04000000 : _GEN_234);
	wire [31:0] _GEN_236 = (10'h0ec == index ? 32'h0f000000 : _GEN_235);
	wire [31:0] _GEN_237 = (10'h0ed == index ? 32'h01000000 : _GEN_236);
	wire [31:0] _GEN_238 = (10'h0ee == index ? 32'h03000000 : _GEN_237);
	wire [31:0] _GEN_239 = (10'h0ef == index ? 32'h2c000000 : _GEN_238);
	wire [31:0] _GEN_240 = (10'h0f0 == index ? 32'h1b000000 : _GEN_239);
	wire [31:0] _GEN_241 = (10'h0f1 == index ? 32'h65657266 : _GEN_240);
	wire [31:0] _GEN_242 = (10'h0f2 == index ? 32'h70696863 : _GEN_241);
	wire [31:0] _GEN_243 = (10'h0f3 == index ? 32'h6f722c73 : _GEN_242);
	wire [31:0] _GEN_244 = (10'h0f4 == index ? 32'h74656b63 : _GEN_243);
	wire [31:0] _GEN_245 = (10'h0f5 == index ? 32'h70696863 : _GEN_244);
	wire [31:0] _GEN_246 = (10'h0f6 == index ? 32'h6b6e752d : _GEN_245);
	wire [31:0] _GEN_247 = (10'h0f7 == index ? 32'h6e776f6e : _GEN_246);
	wire [31:0] _GEN_248 = (10'h0f8 == index ? 32'h636f732d : _GEN_247);
	wire [31:0] _GEN_249 = (10'h0f9 == index ? 32'h6d697300 : _GEN_248);
	wire [31:0] _GEN_250 = (10'h0fa == index ? 32'h2d656c70 : _GEN_249);
	wire [31:0] _GEN_251 = (10'h0fb == index ? 32'h00737562 : _GEN_250);
	wire [31:0] _GEN_252 = (10'h0fc == index ? 32'h03000000 : _GEN_251);
	wire [31:0] _GEN_253 = (10'h0fd == index ? 32'h00000000 : _GEN_252);
	wire [31:0] _GEN_254 = (10'h0fe == index ? 32'h24010000 : _GEN_253);
	wire [31:0] _GEN_255 = (10'h0ff == index ? 32'h01000000 : _GEN_254);
	wire [31:0] _GEN_256 = (10'h100 == index ? 32'h746f6f62 : _GEN_255);
	wire [31:0] _GEN_257 = (10'h101 == index ? 32'h6464612d : _GEN_256);
	wire [31:0] _GEN_258 = (10'h102 == index ? 32'h73736572 : _GEN_257);
	wire [31:0] _GEN_259 = (10'h103 == index ? 32'h6765722d : _GEN_258);
	wire [31:0] _GEN_260 = (10'h104 == index ? 32'h30303440 : _GEN_259);
	wire [31:0] _GEN_261 = (10'h105 == index ? 32'h00000030 : _GEN_260);
	wire [31:0] _GEN_262 = (10'h106 == index ? 32'h03000000 : _GEN_261);
	wire [31:0] _GEN_263 = (10'h107 == index ? 32'h08000000 : _GEN_262);
	wire [31:0] _GEN_264 = (10'h108 == index ? 32'haf000000 : _GEN_263);
	wire [31:0] _GEN_265 = (10'h109 == index ? 32'h00400000 : _GEN_264);
	wire [31:0] _GEN_266 = (10'h10a == index ? 32'h00100000 : _GEN_265);
	wire [31:0] _GEN_267 = (10'h10b == index ? 32'h03000000 : _GEN_266);
	wire [31:0] _GEN_268 = (10'h10c == index ? 32'h08000000 : _GEN_267);
	wire [31:0] _GEN_269 = (10'h10d == index ? 32'h2b010000 : _GEN_268);
	wire [31:0] _GEN_270 = (10'h10e == index ? 32'h746e6f63 : _GEN_269);
	wire [31:0] _GEN_271 = (10'h10f == index ? 32'h006c6f72 : _GEN_270);
	wire [31:0] _GEN_272 = (10'h110 == index ? 32'h02000000 : _GEN_271);
	wire [31:0] _GEN_273 = (10'h111 == index ? 32'h01000000 : _GEN_272);
	wire [31:0] _GEN_274 = (10'h112 == index ? 32'h6e696c63 : _GEN_273);
	wire [31:0] _GEN_275 = (10'h113 == index ? 32'h30324074 : _GEN_274);
	wire [31:0] _GEN_276 = (10'h114 == index ? 32'h30303030 : _GEN_275);
	wire [31:0] _GEN_277 = (10'h115 == index ? 32'h00000030 : _GEN_276);
	wire [31:0] _GEN_278 = (10'h116 == index ? 32'h03000000 : _GEN_277);
	wire [31:0] _GEN_279 = (10'h117 == index ? 32'h0d000000 : _GEN_278);
	wire [31:0] _GEN_280 = (10'h118 == index ? 32'h1b000000 : _GEN_279);
	wire [31:0] _GEN_281 = (10'h119 == index ? 32'h63736972 : _GEN_280);
	wire [31:0] _GEN_282 = (10'h11a == index ? 32'h6c632c76 : _GEN_281);
	wire [31:0] _GEN_283 = (10'h11b == index ? 32'h30746e69 : _GEN_282);
	wire [31:0] _GEN_284 = (10'h11c == index ? 32'h00000000 : _GEN_283);
	wire [31:0] _GEN_285 = (10'h11d == index ? 32'h03000000 : _GEN_284);
	wire [31:0] _GEN_286 = (10'h11e == index ? 32'h10000000 : _GEN_285);
	wire [31:0] _GEN_287 = (10'h11f == index ? 32'h35010000 : _GEN_286);
	wire [31:0] _GEN_288 = (10'h120 == index ? 32'h02000000 : _GEN_287);
	wire [31:0] _GEN_289 = (10'h121 == index ? 32'h03000000 : _GEN_288);
	wire [31:0] _GEN_290 = (10'h122 == index ? 32'h02000000 : _GEN_289);
	wire [31:0] _GEN_291 = (10'h123 == index ? 32'h07000000 : _GEN_290);
	wire [31:0] _GEN_292 = (10'h124 == index ? 32'h03000000 : _GEN_291);
	wire [31:0] _GEN_293 = (10'h125 == index ? 32'h08000000 : _GEN_292);
	wire [31:0] _GEN_294 = (10'h126 == index ? 32'haf000000 : _GEN_293);
	wire [31:0] _GEN_295 = (10'h127 == index ? 32'h00000002 : _GEN_294);
	wire [31:0] _GEN_296 = (10'h128 == index ? 32'h00000100 : _GEN_295);
	wire [31:0] _GEN_297 = (10'h129 == index ? 32'h03000000 : _GEN_296);
	wire [31:0] _GEN_298 = (10'h12a == index ? 32'h08000000 : _GEN_297);
	wire [31:0] _GEN_299 = (10'h12b == index ? 32'h2b010000 : _GEN_298);
	wire [31:0] _GEN_300 = (10'h12c == index ? 32'h746e6f63 : _GEN_299);
	wire [31:0] _GEN_301 = (10'h12d == index ? 32'h006c6f72 : _GEN_300);
	wire [31:0] _GEN_302 = (10'h12e == index ? 32'h02000000 : _GEN_301);
	wire [31:0] _GEN_303 = (10'h12f == index ? 32'h01000000 : _GEN_302);
	wire [31:0] _GEN_304 = (10'h130 == index ? 32'h636f6c63 : _GEN_303);
	wire [31:0] _GEN_305 = (10'h131 == index ? 32'h61672d6b : _GEN_304);
	wire [31:0] _GEN_306 = (10'h132 == index ? 32'h40726574 : _GEN_305);
	wire [31:0] _GEN_307 = (10'h133 == index ? 32'h30303031 : _GEN_306);
	wire [31:0] _GEN_308 = (10'h134 == index ? 32'h00003030 : _GEN_307);
	wire [31:0] _GEN_309 = (10'h135 == index ? 32'h03000000 : _GEN_308);
	wire [31:0] _GEN_310 = (10'h136 == index ? 32'h08000000 : _GEN_309);
	wire [31:0] _GEN_311 = (10'h137 == index ? 32'haf000000 : _GEN_310);
	wire [31:0] _GEN_312 = (10'h138 == index ? 32'h00001000 : _GEN_311);
	wire [31:0] _GEN_313 = (10'h139 == index ? 32'h00100000 : _GEN_312);
	wire [31:0] _GEN_314 = (10'h13a == index ? 32'h03000000 : _GEN_313);
	wire [31:0] _GEN_315 = (10'h13b == index ? 32'h08000000 : _GEN_314);
	wire [31:0] _GEN_316 = (10'h13c == index ? 32'h2b010000 : _GEN_315);
	wire [31:0] _GEN_317 = (10'h13d == index ? 32'h746e6f63 : _GEN_316);
	wire [31:0] _GEN_318 = (10'h13e == index ? 32'h006c6f72 : _GEN_317);
	wire [31:0] _GEN_319 = (10'h13f == index ? 32'h02000000 : _GEN_318);
	wire [31:0] _GEN_320 = (10'h140 == index ? 32'h01000000 : _GEN_319);
	wire [31:0] _GEN_321 = (10'h141 == index ? 32'h75626564 : _GEN_320);
	wire [31:0] _GEN_322 = (10'h142 == index ? 32'h6f632d67 : _GEN_321);
	wire [31:0] _GEN_323 = (10'h143 == index ? 32'h6f72746e : _GEN_322);
	wire [31:0] _GEN_324 = (10'h144 == index ? 32'h72656c6c : _GEN_323);
	wire [31:0] _GEN_325 = (10'h145 == index ? 32'h00003040 : _GEN_324);
	wire [31:0] _GEN_326 = (10'h146 == index ? 32'h03000000 : _GEN_325);
	wire [31:0] _GEN_327 = (10'h147 == index ? 32'h21000000 : _GEN_326);
	wire [31:0] _GEN_328 = (10'h148 == index ? 32'h1b000000 : _GEN_327);
	wire [31:0] _GEN_329 = (10'h149 == index ? 32'h69666973 : _GEN_328);
	wire [31:0] _GEN_330 = (10'h14a == index ? 32'h642c6576 : _GEN_329);
	wire [31:0] _GEN_331 = (10'h14b == index ? 32'h67756265 : _GEN_330);
	wire [31:0] _GEN_332 = (10'h14c == index ? 32'h3331302d : _GEN_331);
	wire [31:0] _GEN_333 = (10'h14d == index ? 32'h73697200 : _GEN_332);
	wire [31:0] _GEN_334 = (10'h14e == index ? 32'h642c7663 : _GEN_333);
	wire [31:0] _GEN_335 = (10'h14f == index ? 32'h67756265 : _GEN_334);
	wire [31:0] _GEN_336 = (10'h150 == index ? 32'h3331302d : _GEN_335);
	wire [31:0] _GEN_337 = (10'h151 == index ? 32'h00000000 : _GEN_336);
	wire [31:0] _GEN_338 = (10'h152 == index ? 32'h03000000 : _GEN_337);
	wire [31:0] _GEN_339 = (10'h153 == index ? 32'h05000000 : _GEN_338);
	wire [31:0] _GEN_340 = (10'h154 == index ? 32'h49010000 : _GEN_339);
	wire [31:0] _GEN_341 = (10'h155 == index ? 32'h6761746a : _GEN_340);
	wire [31:0] _GEN_342 = (10'h156 == index ? 32'h00000000 : _GEN_341);
	wire [31:0] _GEN_343 = (10'h157 == index ? 32'h03000000 : _GEN_342);
	wire [31:0] _GEN_344 = (10'h158 == index ? 32'h08000000 : _GEN_343);
	wire [31:0] _GEN_345 = (10'h159 == index ? 32'h35010000 : _GEN_344);
	wire [31:0] _GEN_346 = (10'h15a == index ? 32'h02000000 : _GEN_345);
	wire [31:0] _GEN_347 = (10'h15b == index ? 32'hffff0000 : _GEN_346);
	wire [31:0] _GEN_348 = (10'h15c == index ? 32'h03000000 : _GEN_347);
	wire [31:0] _GEN_349 = (10'h15d == index ? 32'h08000000 : _GEN_348);
	wire [31:0] _GEN_350 = (10'h15e == index ? 32'haf000000 : _GEN_349);
	wire [31:0] _GEN_351 = (10'h15f == index ? 32'h00000000 : _GEN_350);
	wire [31:0] _GEN_352 = (10'h160 == index ? 32'h00100000 : _GEN_351);
	wire [31:0] _GEN_353 = (10'h161 == index ? 32'h03000000 : _GEN_352);
	wire [31:0] _GEN_354 = (10'h162 == index ? 32'h08000000 : _GEN_353);
	wire [31:0] _GEN_355 = (10'h163 == index ? 32'h2b010000 : _GEN_354);
	wire [31:0] _GEN_356 = (10'h164 == index ? 32'h746e6f63 : _GEN_355);
	wire [31:0] _GEN_357 = (10'h165 == index ? 32'h006c6f72 : _GEN_356);
	wire [31:0] _GEN_358 = (10'h166 == index ? 32'h02000000 : _GEN_357);
	wire [31:0] _GEN_359 = (10'h167 == index ? 32'h01000000 : _GEN_358);
	wire [31:0] _GEN_360 = (10'h168 == index ? 32'h6d697464 : _GEN_359);
	wire [31:0] _GEN_361 = (10'h169 == index ? 32'h30303840 : _GEN_360);
	wire [31:0] _GEN_362 = (10'h16a == index ? 32'h30303030 : _GEN_361);
	wire [31:0] _GEN_363 = (10'h16b == index ? 32'h00000030 : _GEN_362);
	wire [31:0] _GEN_364 = (10'h16c == index ? 32'h03000000 : _GEN_363);
	wire [31:0] _GEN_365 = (10'h16d == index ? 32'h0d000000 : _GEN_364);
	wire [31:0] _GEN_366 = (10'h16e == index ? 32'h1b000000 : _GEN_365);
	wire [31:0] _GEN_367 = (10'h16f == index ? 32'h69666973 : _GEN_366);
	wire [31:0] _GEN_368 = (10'h170 == index ? 32'h642c6576 : _GEN_367);
	wire [31:0] _GEN_369 = (10'h171 == index ? 32'h306d6974 : _GEN_368);
	wire [31:0] _GEN_370 = (10'h172 == index ? 32'h00000000 : _GEN_369);
	wire [31:0] _GEN_371 = (10'h173 == index ? 32'h03000000 : _GEN_370);
	wire [31:0] _GEN_372 = (10'h174 == index ? 32'h08000000 : _GEN_371);
	wire [31:0] _GEN_373 = (10'h175 == index ? 32'haf000000 : _GEN_372);
	wire [31:0] _GEN_374 = (10'h176 == index ? 32'h00000080 : _GEN_373);
	wire [31:0] _GEN_375 = (10'h177 == index ? 32'h00400000 : _GEN_374);
	wire [31:0] _GEN_376 = (10'h178 == index ? 32'h03000000 : _GEN_375);
	wire [31:0] _GEN_377 = (10'h179 == index ? 32'h04000000 : _GEN_376);
	wire [31:0] _GEN_378 = (10'h17a == index ? 32'h2b010000 : _GEN_377);
	wire [31:0] _GEN_379 = (10'h17b == index ? 32'h006d656d : _GEN_378);
	wire [31:0] _GEN_380 = (10'h17c == index ? 32'h03000000 : _GEN_379);
	wire [31:0] _GEN_381 = (10'h17d == index ? 32'h04000000 : _GEN_380);
	wire [31:0] _GEN_382 = (10'h17e == index ? 32'h1c010000 : _GEN_381);
	wire [31:0] _GEN_383 = (10'h17f == index ? 32'h01000000 : _GEN_382);
	wire [31:0] _GEN_384 = (10'h180 == index ? 32'h02000000 : _GEN_383);
	wire [31:0] _GEN_385 = (10'h181 == index ? 32'h01000000 : _GEN_384);
	wire [31:0] _GEN_386 = (10'h182 == index ? 32'h6f727265 : _GEN_385);
	wire [31:0] _GEN_387 = (10'h183 == index ? 32'h65642d72 : _GEN_386);
	wire [31:0] _GEN_388 = (10'h184 == index ? 32'h65636976 : _GEN_387);
	wire [31:0] _GEN_389 = (10'h185 == index ? 32'h30303340 : _GEN_388);
	wire [31:0] _GEN_390 = (10'h186 == index ? 32'h00000030 : _GEN_389);
	wire [31:0] _GEN_391 = (10'h187 == index ? 32'h03000000 : _GEN_390);
	wire [31:0] _GEN_392 = (10'h188 == index ? 32'h0e000000 : _GEN_391);
	wire [31:0] _GEN_393 = (10'h189 == index ? 32'h1b000000 : _GEN_392);
	wire [31:0] _GEN_394 = (10'h18a == index ? 32'h69666973 : _GEN_393);
	wire [31:0] _GEN_395 = (10'h18b == index ? 32'h652c6576 : _GEN_394);
	wire [31:0] _GEN_396 = (10'h18c == index ? 32'h726f7272 : _GEN_395);
	wire [31:0] _GEN_397 = (10'h18d == index ? 32'h00000030 : _GEN_396);
	wire [31:0] _GEN_398 = (10'h18e == index ? 32'h03000000 : _GEN_397);
	wire [31:0] _GEN_399 = (10'h18f == index ? 32'h08000000 : _GEN_398);
	wire [31:0] _GEN_400 = (10'h190 == index ? 32'haf000000 : _GEN_399);
	wire [31:0] _GEN_401 = (10'h191 == index ? 32'h00300000 : _GEN_400);
	wire [31:0] _GEN_402 = (10'h192 == index ? 32'h00100000 : _GEN_401);
	wire [31:0] _GEN_403 = (10'h193 == index ? 32'h02000000 : _GEN_402);
	wire [31:0] _GEN_404 = (10'h194 == index ? 32'h01000000 : _GEN_403);
	wire [31:0] _GEN_405 = (10'h195 == index ? 32'h65746e69 : _GEN_404);
	wire [31:0] _GEN_406 = (10'h196 == index ? 32'h70757272 : _GEN_405);
	wire [31:0] _GEN_407 = (10'h197 == index ? 32'h6f632d74 : _GEN_406);
	wire [31:0] _GEN_408 = (10'h198 == index ? 32'h6f72746e : _GEN_407);
	wire [31:0] _GEN_409 = (10'h199 == index ? 32'h72656c6c : _GEN_408);
	wire [31:0] _GEN_410 = (10'h19a == index ? 32'h30306340 : _GEN_409);
	wire [31:0] _GEN_411 = (10'h19b == index ? 32'h30303030 : _GEN_410);
	wire [31:0] _GEN_412 = (10'h19c == index ? 32'h00000000 : _GEN_411);
	wire [31:0] _GEN_413 = (10'h19d == index ? 32'h03000000 : _GEN_412);
	wire [31:0] _GEN_414 = (10'h19e == index ? 32'h04000000 : _GEN_413);
	wire [31:0] _GEN_415 = (10'h19f == index ? 32'hf6000000 : _GEN_414);
	wire [31:0] _GEN_416 = (10'h1a0 == index ? 32'h01000000 : _GEN_415);
	wire [31:0] _GEN_417 = (10'h1a1 == index ? 32'h03000000 : _GEN_416);
	wire [31:0] _GEN_418 = (10'h1a2 == index ? 32'h0c000000 : _GEN_417);
	wire [31:0] _GEN_419 = (10'h1a3 == index ? 32'h1b000000 : _GEN_418);
	wire [31:0] _GEN_420 = (10'h1a4 == index ? 32'h63736972 : _GEN_419);
	wire [31:0] _GEN_421 = (10'h1a5 == index ? 32'h6c702c76 : _GEN_420);
	wire [31:0] _GEN_422 = (10'h1a6 == index ? 32'h00306369 : _GEN_421);
	wire [31:0] _GEN_423 = (10'h1a7 == index ? 32'h03000000 : _GEN_422);
	wire [31:0] _GEN_424 = (10'h1a8 == index ? 32'h00000000 : _GEN_423);
	wire [31:0] _GEN_425 = (10'h1a9 == index ? 32'h07010000 : _GEN_424);
	wire [31:0] _GEN_426 = (10'h1aa == index ? 32'h03000000 : _GEN_425);
	wire [31:0] _GEN_427 = (10'h1ab == index ? 32'h08000000 : _GEN_426);
	wire [31:0] _GEN_428 = (10'h1ac == index ? 32'h35010000 : _GEN_427);
	wire [31:0] _GEN_429 = (10'h1ad == index ? 32'h02000000 : _GEN_428);
	wire [31:0] _GEN_430 = (10'h1ae == index ? 32'h0b000000 : _GEN_429);
	wire [31:0] _GEN_431 = (10'h1af == index ? 32'h03000000 : _GEN_430);
	wire [31:0] _GEN_432 = (10'h1b0 == index ? 32'h08000000 : _GEN_431);
	wire [31:0] _GEN_433 = (10'h1b1 == index ? 32'haf000000 : _GEN_432);
	wire [31:0] _GEN_434 = (10'h1b2 == index ? 32'h0000000c : _GEN_433);
	wire [31:0] _GEN_435 = (10'h1b3 == index ? 32'h00000004 : _GEN_434);
	wire [31:0] _GEN_436 = (10'h1b4 == index ? 32'h03000000 : _GEN_435);
	wire [31:0] _GEN_437 = (10'h1b5 == index ? 32'h08000000 : _GEN_436);
	wire [31:0] _GEN_438 = (10'h1b6 == index ? 32'h2b010000 : _GEN_437);
	wire [31:0] _GEN_439 = (10'h1b7 == index ? 32'h746e6f63 : _GEN_438);
	wire [31:0] _GEN_440 = (10'h1b8 == index ? 32'h006c6f72 : _GEN_439);
	wire [31:0] _GEN_441 = (10'h1b9 == index ? 32'h03000000 : _GEN_440);
	wire [31:0] _GEN_442 = (10'h1ba == index ? 32'h04000000 : _GEN_441);
	wire [31:0] _GEN_443 = (10'h1bb == index ? 32'h56010000 : _GEN_442);
	wire [31:0] _GEN_444 = (10'h1bc == index ? 32'h01000000 : _GEN_443);
	wire [31:0] _GEN_445 = (10'h1bd == index ? 32'h03000000 : _GEN_444);
	wire [31:0] _GEN_446 = (10'h1be == index ? 32'h04000000 : _GEN_445);
	wire [31:0] _GEN_447 = (10'h1bf == index ? 32'h69010000 : _GEN_446);
	wire [31:0] _GEN_448 = (10'h1c0 == index ? 32'h01000000 : _GEN_447);
	wire [31:0] _GEN_449 = (10'h1c1 == index ? 32'h03000000 : _GEN_448);
	wire [31:0] _GEN_450 = (10'h1c2 == index ? 32'h04000000 : _GEN_449);
	wire [31:0] _GEN_451 = (10'h1c3 == index ? 32'h1c010000 : _GEN_450);
	wire [31:0] _GEN_452 = (10'h1c4 == index ? 32'h04000000 : _GEN_451);
	wire [31:0] _GEN_453 = (10'h1c5 == index ? 32'h02000000 : _GEN_452);
	wire [31:0] _GEN_454 = (10'h1c6 == index ? 32'h01000000 : _GEN_453);
	wire [31:0] _GEN_455 = (10'h1c7 == index ? 32'h6977626c : _GEN_454);
	wire [31:0] _GEN_456 = (10'h1c8 == index ? 32'h61722d66 : _GEN_455);
	wire [31:0] _GEN_457 = (10'h1c9 == index ? 32'h3031406d : _GEN_456);
	wire [31:0] _GEN_458 = (10'h1ca == index ? 32'h30303030 : _GEN_457);
	wire [31:0] _GEN_459 = (10'h1cb == index ? 32'h00003030 : _GEN_458);
	wire [31:0] _GEN_460 = (10'h1cc == index ? 32'h03000000 : _GEN_459);
	wire [31:0] _GEN_461 = (10'h1cd == index ? 32'h08000000 : _GEN_460);
	wire [31:0] _GEN_462 = (10'h1ce == index ? 32'haf000000 : _GEN_461);
	wire [31:0] _GEN_463 = (10'h1cf == index ? 32'h00000010 : _GEN_462);
	wire [31:0] _GEN_464 = (10'h1d0 == index ? 32'h00100000 : _GEN_463);
	wire [31:0] _GEN_465 = (10'h1d1 == index ? 32'h02000000 : _GEN_464);
	wire [31:0] _GEN_466 = (10'h1d2 == index ? 32'h01000000 : _GEN_465);
	wire [31:0] _GEN_467 = (10'h1d3 == index ? 32'h6977626c : _GEN_466);
	wire [31:0] _GEN_468 = (10'h1d4 == index ? 32'h6f722d66 : _GEN_467);
	wire [31:0] _GEN_469 = (10'h1d5 == index ? 32'h3032406d : _GEN_468);
	wire [31:0] _GEN_470 = (10'h1d6 == index ? 32'h00303030 : _GEN_469);
	wire [31:0] _GEN_471 = (10'h1d7 == index ? 32'h03000000 : _GEN_470);
	wire [31:0] _GEN_472 = (10'h1d8 == index ? 32'h08000000 : _GEN_471);
	wire [31:0] _GEN_473 = (10'h1d9 == index ? 32'haf000000 : _GEN_472);
	wire [31:0] _GEN_474 = (10'h1da == index ? 32'h00000200 : _GEN_473);
	wire [31:0] _GEN_475 = (10'h1db == index ? 32'h00000100 : _GEN_474);
	wire [31:0] _GEN_476 = (10'h1dc == index ? 32'h02000000 : _GEN_475);
	wire [31:0] _GEN_477 = (10'h1dd == index ? 32'h01000000 : _GEN_476);
	wire [31:0] _GEN_478 = (10'h1de == index ? 32'h406d6f72 : _GEN_477);
	wire [31:0] _GEN_479 = (10'h1df == index ? 32'h30303031 : _GEN_478);
	wire [31:0] _GEN_480 = (10'h1e0 == index ? 32'h00000030 : _GEN_479);
	wire [31:0] _GEN_481 = (10'h1e1 == index ? 32'h03000000 : _GEN_480);
	wire [31:0] _GEN_482 = (10'h1e2 == index ? 32'h0c000000 : _GEN_481);
	wire [31:0] _GEN_483 = (10'h1e3 == index ? 32'h1b000000 : _GEN_482);
	wire [31:0] _GEN_484 = (10'h1e4 == index ? 32'h69666973 : _GEN_483);
	wire [31:0] _GEN_485 = (10'h1e5 == index ? 32'h722c6576 : _GEN_484);
	wire [31:0] _GEN_486 = (10'h1e6 == index ? 32'h00306d6f : _GEN_485);
	wire [31:0] _GEN_487 = (10'h1e7 == index ? 32'h03000000 : _GEN_486);
	wire [31:0] _GEN_488 = (10'h1e8 == index ? 32'h08000000 : _GEN_487);
	wire [31:0] _GEN_489 = (10'h1e9 == index ? 32'haf000000 : _GEN_488);
	wire [31:0] _GEN_490 = (10'h1ea == index ? 32'h00000100 : _GEN_489);
	wire [31:0] _GEN_491 = (10'h1eb == index ? 32'h00000100 : _GEN_490);
	wire [31:0] _GEN_492 = (10'h1ec == index ? 32'h03000000 : _GEN_491);
	wire [31:0] _GEN_493 = (10'h1ed == index ? 32'h04000000 : _GEN_492);
	wire [31:0] _GEN_494 = (10'h1ee == index ? 32'h2b010000 : _GEN_493);
	wire [31:0] _GEN_495 = (10'h1ef == index ? 32'h006d656d : _GEN_494);
	wire [31:0] _GEN_496 = (10'h1f0 == index ? 32'h02000000 : _GEN_495);
	wire [31:0] _GEN_497 = (10'h1f1 == index ? 32'h01000000 : _GEN_496);
	wire [31:0] _GEN_498 = (10'h1f2 == index ? 32'h69726573 : _GEN_497);
	wire [31:0] _GEN_499 = (10'h1f3 == index ? 32'h35406c61 : _GEN_498);
	wire [31:0] _GEN_500 = (10'h1f4 == index ? 32'h30303034 : _GEN_499);
	wire [31:0] _GEN_501 = (10'h1f5 == index ? 32'h00303030 : _GEN_500);
	wire [31:0] _GEN_502 = (10'h1f6 == index ? 32'h03000000 : _GEN_501);
	wire [31:0] _GEN_503 = (10'h1f7 == index ? 32'h04000000 : _GEN_502);
	wire [31:0] _GEN_504 = (10'h1f8 == index ? 32'h74010000 : _GEN_503);
	wire [31:0] _GEN_505 = (10'h1f9 == index ? 32'h03000000 : _GEN_504);
	wire [31:0] _GEN_506 = (10'h1fa == index ? 32'h03000000 : _GEN_505);
	wire [31:0] _GEN_507 = (10'h1fb == index ? 32'h0d000000 : _GEN_506);
	wire [31:0] _GEN_508 = (10'h1fc == index ? 32'h1b000000 : _GEN_507);
	wire [31:0] _GEN_509 = (10'h1fd == index ? 32'h69666973 : _GEN_508);
	wire [31:0] _GEN_510 = (10'h1fe == index ? 32'h752c6576 : _GEN_509);
	wire [31:0] _GEN_511 = (10'h1ff == index ? 32'h30747261 : _GEN_510);
	wire [31:0] _GEN_512 = (10'h200 == index ? 32'h00000000 : _GEN_511);
	wire [31:0] _GEN_513 = (10'h201 == index ? 32'h03000000 : _GEN_512);
	wire [31:0] _GEN_514 = (10'h202 == index ? 32'h04000000 : _GEN_513);
	wire [31:0] _GEN_515 = (10'h203 == index ? 32'h7b010000 : _GEN_514);
	wire [31:0] _GEN_516 = (10'h204 == index ? 32'h04000000 : _GEN_515);
	wire [31:0] _GEN_517 = (10'h205 == index ? 32'h03000000 : _GEN_516);
	wire [31:0] _GEN_518 = (10'h206 == index ? 32'h04000000 : _GEN_517);
	wire [31:0] _GEN_519 = (10'h207 == index ? 32'h8c010000 : _GEN_518);
	wire [31:0] _GEN_520 = (10'h208 == index ? 32'h01000000 : _GEN_519);
	wire [31:0] _GEN_521 = (10'h209 == index ? 32'h03000000 : _GEN_520);
	wire [31:0] _GEN_522 = (10'h20a == index ? 32'h08000000 : _GEN_521);
	wire [31:0] _GEN_523 = (10'h20b == index ? 32'haf000000 : _GEN_522);
	wire [31:0] _GEN_524 = (10'h20c == index ? 32'h00000054 : _GEN_523);
	wire [31:0] _GEN_525 = (10'h20d == index ? 32'h00100000 : _GEN_524);
	wire [31:0] _GEN_526 = (10'h20e == index ? 32'h03000000 : _GEN_525);
	wire [31:0] _GEN_527 = (10'h20f == index ? 32'h08000000 : _GEN_526);
	wire [31:0] _GEN_528 = (10'h210 == index ? 32'h2b010000 : _GEN_527);
	wire [31:0] _GEN_529 = (10'h211 == index ? 32'h746e6f63 : _GEN_528);
	wire [31:0] _GEN_530 = (10'h212 == index ? 32'h006c6f72 : _GEN_529);
	wire [31:0] _GEN_531 = (10'h213 == index ? 32'h02000000 : _GEN_530);
	wire [31:0] _GEN_532 = (10'h214 == index ? 32'h01000000 : _GEN_531);
	wire [31:0] _GEN_533 = (10'h215 == index ? 32'h73627573 : _GEN_532);
	wire [31:0] _GEN_534 = (10'h216 == index ? 32'h65747379 : _GEN_533);
	wire [31:0] _GEN_535 = (10'h217 == index ? 32'h62705f6d : _GEN_534);
	wire [31:0] _GEN_536 = (10'h218 == index ? 32'h635f7375 : _GEN_535);
	wire [31:0] _GEN_537 = (10'h219 == index ? 32'h6b636f6c : _GEN_536);
	wire [31:0] _GEN_538 = (10'h21a == index ? 32'h00000000 : _GEN_537);
	wire [31:0] _GEN_539 = (10'h21b == index ? 32'h03000000 : _GEN_538);
	wire [31:0] _GEN_540 = (10'h21c == index ? 32'h04000000 : _GEN_539);
	wire [31:0] _GEN_541 = (10'h21d == index ? 32'h97010000 : _GEN_540);
	wire [31:0] _GEN_542 = (10'h21e == index ? 32'h00000000 : _GEN_541);
	wire [31:0] _GEN_543 = (10'h21f == index ? 32'h03000000 : _GEN_542);
	wire [31:0] _GEN_544 = (10'h220 == index ? 32'h04000000 : _GEN_543);
	wire [31:0] _GEN_545 = (10'h221 == index ? 32'h47000000 : _GEN_544);
	wire [31:0] _GEN_546 = (10'h222 == index ? 32'h00e1f505 : _GEN_545);
	wire [31:0] _GEN_547 = (10'h223 == index ? 32'h03000000 : _GEN_546);
	wire [31:0] _GEN_548 = (10'h224 == index ? 32'h15000000 : _GEN_547);
	wire [31:0] _GEN_549 = (10'h225 == index ? 32'ha4010000 : _GEN_548);
	wire [31:0] _GEN_550 = (10'h226 == index ? 32'h73627573 : _GEN_549);
	wire [31:0] _GEN_551 = (10'h227 == index ? 32'h65747379 : _GEN_550);
	wire [31:0] _GEN_552 = (10'h228 == index ? 32'h62705f6d : _GEN_551);
	wire [31:0] _GEN_553 = (10'h229 == index ? 32'h635f7375 : _GEN_552);
	wire [31:0] _GEN_554 = (10'h22a == index ? 32'h6b636f6c : _GEN_553);
	wire [31:0] _GEN_555 = (10'h22b == index ? 32'h00000000 : _GEN_554);
	wire [31:0] _GEN_556 = (10'h22c == index ? 32'h03000000 : _GEN_555);
	wire [31:0] _GEN_557 = (10'h22d == index ? 32'h0c000000 : _GEN_556);
	wire [31:0] _GEN_558 = (10'h22e == index ? 32'h1b000000 : _GEN_557);
	wire [31:0] _GEN_559 = (10'h22f == index ? 32'h65786966 : _GEN_558);
	wire [31:0] _GEN_560 = (10'h230 == index ? 32'h6c632d64 : _GEN_559);
	wire [31:0] _GEN_561 = (10'h231 == index ? 32'h006b636f : _GEN_560);
	wire [31:0] _GEN_562 = (10'h232 == index ? 32'h03000000 : _GEN_561);
	wire [31:0] _GEN_563 = (10'h233 == index ? 32'h04000000 : _GEN_562);
	wire [31:0] _GEN_564 = (10'h234 == index ? 32'h1c010000 : _GEN_563);
	wire [31:0] _GEN_565 = (10'h235 == index ? 32'h03000000 : _GEN_564);
	wire [31:0] _GEN_566 = (10'h236 == index ? 32'h02000000 : _GEN_565);
	wire [31:0] _GEN_567 = (10'h237 == index ? 32'h01000000 : _GEN_566);
	wire [31:0] _GEN_568 = (10'h238 == index ? 32'h656c6974 : _GEN_567);
	wire [31:0] _GEN_569 = (10'h239 == index ? 32'h7365722d : _GEN_568);
	wire [31:0] _GEN_570 = (10'h23a == index ? 32'h732d7465 : _GEN_569);
	wire [31:0] _GEN_571 = (10'h23b == index ? 32'h65747465 : _GEN_570);
	wire [31:0] _GEN_572 = (10'h23c == index ? 32'h31314072 : _GEN_571);
	wire [31:0] _GEN_573 = (10'h23d == index ? 32'h30303030 : _GEN_572);
	wire [31:0] _GEN_574 = (10'h23e == index ? 32'h00000000 : _GEN_573);
	wire [31:0] _GEN_575 = (10'h23f == index ? 32'h03000000 : _GEN_574);
	wire [31:0] _GEN_576 = (10'h240 == index ? 32'h08000000 : _GEN_575);
	wire [31:0] _GEN_577 = (10'h241 == index ? 32'haf000000 : _GEN_576);
	wire [31:0] _GEN_578 = (10'h242 == index ? 32'h00001100 : _GEN_577);
	wire [31:0] _GEN_579 = (10'h243 == index ? 32'h00100000 : _GEN_578);
	wire [31:0] _GEN_580 = (10'h244 == index ? 32'h03000000 : _GEN_579);
	wire [31:0] _GEN_581 = (10'h245 == index ? 32'h08000000 : _GEN_580);
	wire [31:0] _GEN_582 = (10'h246 == index ? 32'h2b010000 : _GEN_581);
	wire [31:0] _GEN_583 = (10'h247 == index ? 32'h746e6f63 : _GEN_582);
	wire [31:0] _GEN_584 = (10'h248 == index ? 32'h006c6f72 : _GEN_583);
	wire [31:0] _GEN_585 = (10'h249 == index ? 32'h02000000 : _GEN_584);
	wire [31:0] _GEN_586 = (10'h24a == index ? 32'h02000000 : _GEN_585);
	wire [31:0] _GEN_587 = (10'h24b == index ? 32'h02000000 : _GEN_586);
	wire [31:0] _GEN_588 = (10'h24c == index ? 32'h09000000 : _GEN_587);
	wire [31:0] _GEN_589 = (10'h24d == index ? 32'h64646123 : _GEN_588);
	wire [31:0] _GEN_590 = (10'h24e == index ? 32'h73736572 : _GEN_589);
	wire [31:0] _GEN_591 = (10'h24f == index ? 32'h6c65632d : _GEN_590);
	wire [31:0] _GEN_592 = (10'h250 == index ? 32'h2300736c : _GEN_591);
	wire [31:0] _GEN_593 = (10'h251 == index ? 32'h657a6973 : _GEN_592);
	wire [31:0] _GEN_594 = (10'h252 == index ? 32'h6c65632d : _GEN_593);
	wire [31:0] _GEN_595 = (10'h253 == index ? 32'h6300736c : _GEN_594);
	wire [31:0] _GEN_596 = (10'h254 == index ? 32'h61706d6f : _GEN_595);
	wire [31:0] _GEN_597 = (10'h255 == index ? 32'h6c626974 : _GEN_596);
	wire [31:0] _GEN_598 = (10'h256 == index ? 32'h6f6d0065 : _GEN_597);
	wire [31:0] _GEN_599 = (10'h257 == index ? 32'h006c6564 : _GEN_598);
	wire [31:0] _GEN_600 = (10'h258 == index ? 32'h69726573 : _GEN_599);
	wire [31:0] _GEN_601 = (10'h259 == index ? 32'h00306c61 : _GEN_600);
	wire [31:0] _GEN_602 = (10'h25a == index ? 32'h656d6974 : _GEN_601);
	wire [31:0] _GEN_603 = (10'h25b == index ? 32'h65736162 : _GEN_602);
	wire [31:0] _GEN_604 = (10'h25c == index ? 32'h6572662d : _GEN_603);
	wire [31:0] _GEN_605 = (10'h25d == index ? 32'h6e657571 : _GEN_604);
	wire [31:0] _GEN_606 = (10'h25e == index ? 32'h63007963 : _GEN_605);
	wire [31:0] _GEN_607 = (10'h25f == index ? 32'h6b636f6c : _GEN_606);
	wire [31:0] _GEN_608 = (10'h260 == index ? 32'h6572662d : _GEN_607);
	wire [31:0] _GEN_609 = (10'h261 == index ? 32'h6e657571 : _GEN_608);
	wire [31:0] _GEN_610 = (10'h262 == index ? 32'h64007963 : _GEN_609);
	wire [31:0] _GEN_611 = (10'h263 == index ? 32'h63697665 : _GEN_610);
	wire [31:0] _GEN_612 = (10'h264 == index ? 32'h79745f65 : _GEN_611);
	wire [31:0] _GEN_613 = (10'h265 == index ? 32'h68006570 : _GEN_612);
	wire [31:0] _GEN_614 = (10'h266 == index ? 32'h77647261 : _GEN_613);
	wire [31:0] _GEN_615 = (10'h267 == index ? 32'h2d657261 : _GEN_614);
	wire [31:0] _GEN_616 = (10'h268 == index ? 32'h63657865 : _GEN_615);
	wire [31:0] _GEN_617 = (10'h269 == index ? 32'h6572622d : _GEN_616);
	wire [31:0] _GEN_618 = (10'h26a == index ? 32'h6f706b61 : _GEN_617);
	wire [31:0] _GEN_619 = (10'h26b == index ? 32'h2d746e69 : _GEN_618);
	wire [31:0] _GEN_620 = (10'h26c == index ? 32'h6e756f63 : _GEN_619);
	wire [31:0] _GEN_621 = (10'h26d == index ? 32'h2d690074 : _GEN_620);
	wire [31:0] _GEN_622 = (10'h26e == index ? 32'h68636163 : _GEN_621);
	wire [31:0] _GEN_623 = (10'h26f == index ? 32'h6c622d65 : _GEN_622);
	wire [31:0] _GEN_624 = (10'h270 == index ? 32'h2d6b636f : _GEN_623);
	wire [31:0] _GEN_625 = (10'h271 == index ? 32'h657a6973 : _GEN_624);
	wire [31:0] _GEN_626 = (10'h272 == index ? 32'h632d6900 : _GEN_625);
	wire [31:0] _GEN_627 = (10'h273 == index ? 32'h65686361 : _GEN_626);
	wire [31:0] _GEN_628 = (10'h274 == index ? 32'h7465732d : _GEN_627);
	wire [31:0] _GEN_629 = (10'h275 == index ? 32'h2d690073 : _GEN_628);
	wire [31:0] _GEN_630 = (10'h276 == index ? 32'h68636163 : _GEN_629);
	wire [31:0] _GEN_631 = (10'h277 == index ? 32'h69732d65 : _GEN_630);
	wire [31:0] _GEN_632 = (10'h278 == index ? 32'h7200657a : _GEN_631);
	wire [31:0] _GEN_633 = (10'h279 == index ? 32'h72006765 : _GEN_632);
	wire [31:0] _GEN_634 = (10'h27a == index ? 32'h76637369 : _GEN_633);
	wire [31:0] _GEN_635 = (10'h27b == index ? 32'h6173692c : _GEN_634);
	wire [31:0] _GEN_636 = (10'h27c == index ? 32'h73697200 : _GEN_635);
	wire [31:0] _GEN_637 = (10'h27d == index ? 32'h702c7663 : _GEN_636);
	wire [31:0] _GEN_638 = (10'h27e == index ? 32'h7267706d : _GEN_637);
	wire [31:0] _GEN_639 = (10'h27f == index ? 32'h6c756e61 : _GEN_638);
	wire [31:0] _GEN_640 = (10'h280 == index ? 32'h74697261 : _GEN_639);
	wire [31:0] _GEN_641 = (10'h281 == index ? 32'h69720079 : _GEN_640);
	wire [31:0] _GEN_642 = (10'h282 == index ? 32'h2c766373 : _GEN_641);
	wire [31:0] _GEN_643 = (10'h283 == index ? 32'h72706d70 : _GEN_642);
	wire [31:0] _GEN_644 = (10'h284 == index ? 32'h6f696765 : _GEN_643);
	wire [31:0] _GEN_645 = (10'h285 == index ? 32'h7300736e : _GEN_644);
	wire [31:0] _GEN_646 = (10'h286 == index ? 32'h76696669 : _GEN_645);
	wire [31:0] _GEN_647 = (10'h287 == index ? 32'h74642c65 : _GEN_646);
	wire [31:0] _GEN_648 = (10'h288 == index ? 32'h73006d69 : _GEN_647);
	wire [31:0] _GEN_649 = (10'h289 == index ? 32'h75746174 : _GEN_648);
	wire [31:0] _GEN_650 = (10'h28a == index ? 32'h69230073 : _GEN_649);
	wire [31:0] _GEN_651 = (10'h28b == index ? 32'h7265746e : _GEN_650);
	wire [31:0] _GEN_652 = (10'h28c == index ? 32'h74707572 : _GEN_651);
	wire [31:0] _GEN_653 = (10'h28d == index ? 32'h6c65632d : _GEN_652);
	wire [31:0] _GEN_654 = (10'h28e == index ? 32'h6900736c : _GEN_653);
	wire [31:0] _GEN_655 = (10'h28f == index ? 32'h7265746e : _GEN_654);
	wire [31:0] _GEN_656 = (10'h290 == index ? 32'h74707572 : _GEN_655);
	wire [31:0] _GEN_657 = (10'h291 == index ? 32'h6e6f632d : _GEN_656);
	wire [31:0] _GEN_658 = (10'h292 == index ? 32'h6c6f7274 : _GEN_657);
	wire [31:0] _GEN_659 = (10'h293 == index ? 32'h0072656c : _GEN_658);
	wire [31:0] _GEN_660 = (10'h294 == index ? 32'h6e616870 : _GEN_659);
	wire [31:0] _GEN_661 = (10'h295 == index ? 32'h00656c64 : _GEN_660);
	wire [31:0] _GEN_662 = (10'h296 == index ? 32'h676e6172 : _GEN_661);
	wire [31:0] _GEN_663 = (10'h297 == index ? 32'h72007365 : _GEN_662);
	wire [31:0] _GEN_664 = (10'h298 == index ? 32'h6e2d6765 : _GEN_663);
	wire [31:0] _GEN_665 = (10'h299 == index ? 32'h73656d61 : _GEN_664);
	wire [31:0] _GEN_666 = (10'h29a == index ? 32'h746e6900 : _GEN_665);
	wire [31:0] _GEN_667 = (10'h29b == index ? 32'h75727265 : _GEN_666);
	wire [31:0] _GEN_668 = (10'h29c == index ? 32'h2d737470 : _GEN_667);
	wire [31:0] _GEN_669 = (10'h29d == index ? 32'h65747865 : _GEN_668);
	wire [31:0] _GEN_670 = (10'h29e == index ? 32'h6465646e : _GEN_669);
	wire [31:0] _GEN_671 = (10'h29f == index ? 32'h62656400 : _GEN_670);
	wire [31:0] _GEN_672 = (10'h2a0 == index ? 32'h612d6775 : _GEN_671);
	wire [31:0] _GEN_673 = (10'h2a1 == index ? 32'h63617474 : _GEN_672);
	wire [31:0] _GEN_674 = (10'h2a2 == index ? 32'h69720068 : _GEN_673);
	wire [31:0] _GEN_675 = (10'h2a3 == index ? 32'h2c766373 : _GEN_674);
	wire [31:0] _GEN_676 = (10'h2a4 == index ? 32'h2d78616d : _GEN_675);
	wire [31:0] _GEN_677 = (10'h2a5 == index ? 32'h6f697270 : _GEN_676);
	wire [31:0] _GEN_678 = (10'h2a6 == index ? 32'h79746972 : _GEN_677);
	wire [31:0] _GEN_679 = (10'h2a7 == index ? 32'h73697200 : _GEN_678);
	wire [31:0] _GEN_680 = (10'h2a8 == index ? 32'h6e2c7663 : _GEN_679);
	wire [31:0] _GEN_681 = (10'h2a9 == index ? 32'h00766564 : _GEN_680);
	wire [31:0] _GEN_682 = (10'h2aa == index ? 32'h636f6c63 : _GEN_681);
	wire [31:0] _GEN_683 = (10'h2ab == index ? 32'h6900736b : _GEN_682);
	wire [31:0] _GEN_684 = (10'h2ac == index ? 32'h7265746e : _GEN_683);
	wire [31:0] _GEN_685 = (10'h2ad == index ? 32'h74707572 : _GEN_684);
	wire [31:0] _GEN_686 = (10'h2ae == index ? 32'h7261702d : _GEN_685);
	wire [31:0] _GEN_687 = (10'h2af == index ? 32'h00746e65 : _GEN_686);
	wire [31:0] _GEN_688 = (10'h2b0 == index ? 32'h65746e69 : _GEN_687);
	wire [31:0] _GEN_689 = (10'h2b1 == index ? 32'h70757272 : _GEN_688);
	wire [31:0] _GEN_690 = (10'h2b2 == index ? 32'h23007374 : _GEN_689);
	wire [31:0] _GEN_691 = (10'h2b3 == index ? 32'h636f6c63 : _GEN_690);
	wire [31:0] _GEN_692 = (10'h2b4 == index ? 32'h65632d6b : _GEN_691);
	wire [31:0] _GEN_693 = (10'h2b5 == index ? 32'h00736c6c : _GEN_692);
	wire [31:0] _GEN_694 = (10'h2b6 == index ? 32'h636f6c63 : _GEN_693);
	wire [31:0] _GEN_695 = (10'h2b7 == index ? 32'h756f2d6b : _GEN_694);
	wire [31:0] _GEN_696 = (10'h2b8 == index ? 32'h74757074 : _GEN_695);
	wire [31:0] _GEN_697 = (10'h2b9 == index ? 32'h6d616e2d : _GEN_696);
	wire [31:0] _GEN_698 = (10'h2ba == index ? 32'h00007365 : _GEN_697);
	wire [31:0] _GEN_699 = (10'h2bb == index ? 32'h00000000 : _GEN_698);
	wire [31:0] _GEN_700 = (10'h2bc == index ? 32'h00000000 : _GEN_699);
	wire [31:0] _GEN_701 = (10'h2bd == index ? 32'h00000000 : _GEN_700);
	wire [31:0] _GEN_702 = (10'h2be == index ? 32'h00000000 : _GEN_701);
	wire [31:0] _GEN_703 = (10'h2bf == index ? 32'h00000000 : _GEN_702);
	wire [31:0] _GEN_704 = (10'h2c0 == index ? 32'h00000000 : _GEN_703);
	wire [31:0] _GEN_705 = (10'h2c1 == index ? 32'h00000000 : _GEN_704);
	wire [31:0] _GEN_706 = (10'h2c2 == index ? 32'h00000000 : _GEN_705);
	wire [31:0] _GEN_707 = (10'h2c3 == index ? 32'h00000000 : _GEN_706);
	wire [31:0] _GEN_708 = (10'h2c4 == index ? 32'h00000000 : _GEN_707);
	wire [31:0] _GEN_709 = (10'h2c5 == index ? 32'h00000000 : _GEN_708);
	wire [31:0] _GEN_710 = (10'h2c6 == index ? 32'h00000000 : _GEN_709);
	wire [31:0] _GEN_711 = (10'h2c7 == index ? 32'h00000000 : _GEN_710);
	wire [31:0] _GEN_712 = (10'h2c8 == index ? 32'h00000000 : _GEN_711);
	wire [31:0] _GEN_713 = (10'h2c9 == index ? 32'h00000000 : _GEN_712);
	wire [31:0] _GEN_714 = (10'h2ca == index ? 32'h00000000 : _GEN_713);
	wire [31:0] _GEN_715 = (10'h2cb == index ? 32'h00000000 : _GEN_714);
	wire [31:0] _GEN_716 = (10'h2cc == index ? 32'h00000000 : _GEN_715);
	wire [31:0] _GEN_717 = (10'h2cd == index ? 32'h00000000 : _GEN_716);
	wire [31:0] _GEN_718 = (10'h2ce == index ? 32'h00000000 : _GEN_717);
	wire [31:0] _GEN_719 = (10'h2cf == index ? 32'h00000000 : _GEN_718);
	wire [31:0] _GEN_720 = (10'h2d0 == index ? 32'h00000000 : _GEN_719);
	wire [31:0] _GEN_721 = (10'h2d1 == index ? 32'h00000000 : _GEN_720);
	wire [31:0] _GEN_722 = (10'h2d2 == index ? 32'h00000000 : _GEN_721);
	wire [31:0] _GEN_723 = (10'h2d3 == index ? 32'h00000000 : _GEN_722);
	wire [31:0] _GEN_724 = (10'h2d4 == index ? 32'h00000000 : _GEN_723);
	wire [31:0] _GEN_725 = (10'h2d5 == index ? 32'h00000000 : _GEN_724);
	wire [31:0] _GEN_726 = (10'h2d6 == index ? 32'h00000000 : _GEN_725);
	wire [31:0] _GEN_727 = (10'h2d7 == index ? 32'h00000000 : _GEN_726);
	wire [31:0] _GEN_728 = (10'h2d8 == index ? 32'h00000000 : _GEN_727);
	wire [31:0] _GEN_729 = (10'h2d9 == index ? 32'h00000000 : _GEN_728);
	wire [31:0] _GEN_730 = (10'h2da == index ? 32'h00000000 : _GEN_729);
	wire [31:0] _GEN_731 = (10'h2db == index ? 32'h00000000 : _GEN_730);
	wire [31:0] _GEN_732 = (10'h2dc == index ? 32'h00000000 : _GEN_731);
	wire [31:0] _GEN_733 = (10'h2dd == index ? 32'h00000000 : _GEN_732);
	wire [31:0] _GEN_734 = (10'h2de == index ? 32'h00000000 : _GEN_733);
	wire [31:0] _GEN_735 = (10'h2df == index ? 32'h00000000 : _GEN_734);
	wire [31:0] _GEN_736 = (10'h2e0 == index ? 32'h00000000 : _GEN_735);
	wire [31:0] _GEN_737 = (10'h2e1 == index ? 32'h00000000 : _GEN_736);
	wire [31:0] _GEN_738 = (10'h2e2 == index ? 32'h00000000 : _GEN_737);
	wire [31:0] _GEN_739 = (10'h2e3 == index ? 32'h00000000 : _GEN_738);
	wire [31:0] _GEN_740 = (10'h2e4 == index ? 32'h00000000 : _GEN_739);
	wire [31:0] _GEN_741 = (10'h2e5 == index ? 32'h00000000 : _GEN_740);
	wire [31:0] _GEN_742 = (10'h2e6 == index ? 32'h00000000 : _GEN_741);
	wire [31:0] _GEN_743 = (10'h2e7 == index ? 32'h00000000 : _GEN_742);
	wire [31:0] _GEN_744 = (10'h2e8 == index ? 32'h00000000 : _GEN_743);
	wire [31:0] _GEN_745 = (10'h2e9 == index ? 32'h00000000 : _GEN_744);
	wire [31:0] _GEN_746 = (10'h2ea == index ? 32'h00000000 : _GEN_745);
	wire [31:0] _GEN_747 = (10'h2eb == index ? 32'h00000000 : _GEN_746);
	wire [31:0] _GEN_748 = (10'h2ec == index ? 32'h00000000 : _GEN_747);
	wire [31:0] _GEN_749 = (10'h2ed == index ? 32'h00000000 : _GEN_748);
	wire [31:0] _GEN_750 = (10'h2ee == index ? 32'h00000000 : _GEN_749);
	wire [31:0] _GEN_751 = (10'h2ef == index ? 32'h00000000 : _GEN_750);
	wire [31:0] _GEN_752 = (10'h2f0 == index ? 32'h00000000 : _GEN_751);
	wire [31:0] _GEN_753 = (10'h2f1 == index ? 32'h00000000 : _GEN_752);
	wire [31:0] _GEN_754 = (10'h2f2 == index ? 32'h00000000 : _GEN_753);
	wire [31:0] _GEN_755 = (10'h2f3 == index ? 32'h00000000 : _GEN_754);
	wire [31:0] _GEN_756 = (10'h2f4 == index ? 32'h00000000 : _GEN_755);
	wire [31:0] _GEN_757 = (10'h2f5 == index ? 32'h00000000 : _GEN_756);
	wire [31:0] _GEN_758 = (10'h2f6 == index ? 32'h00000000 : _GEN_757);
	wire [31:0] _GEN_759 = (10'h2f7 == index ? 32'h00000000 : _GEN_758);
	wire [31:0] _GEN_760 = (10'h2f8 == index ? 32'h00000000 : _GEN_759);
	wire [31:0] _GEN_761 = (10'h2f9 == index ? 32'h00000000 : _GEN_760);
	wire [31:0] _GEN_762 = (10'h2fa == index ? 32'h00000000 : _GEN_761);
	wire [31:0] _GEN_763 = (10'h2fb == index ? 32'h00000000 : _GEN_762);
	wire [31:0] _GEN_764 = (10'h2fc == index ? 32'h00000000 : _GEN_763);
	wire [31:0] _GEN_765 = (10'h2fd == index ? 32'h00000000 : _GEN_764);
	wire [31:0] _GEN_766 = (10'h2fe == index ? 32'h00000000 : _GEN_765);
	wire [31:0] _GEN_767 = (10'h2ff == index ? 32'h00000000 : _GEN_766);
	wire [31:0] _GEN_768 = (10'h300 == index ? 32'h00000000 : _GEN_767);
	wire [31:0] _GEN_769 = (10'h301 == index ? 32'h00000000 : _GEN_768);
	wire [31:0] _GEN_770 = (10'h302 == index ? 32'h00000000 : _GEN_769);
	wire [31:0] _GEN_771 = (10'h303 == index ? 32'h00000000 : _GEN_770);
	wire [31:0] _GEN_772 = (10'h304 == index ? 32'h00000000 : _GEN_771);
	wire [31:0] _GEN_773 = (10'h305 == index ? 32'h00000000 : _GEN_772);
	wire [31:0] _GEN_774 = (10'h306 == index ? 32'h00000000 : _GEN_773);
	wire [31:0] _GEN_775 = (10'h307 == index ? 32'h00000000 : _GEN_774);
	wire [31:0] _GEN_776 = (10'h308 == index ? 32'h00000000 : _GEN_775);
	wire [31:0] _GEN_777 = (10'h309 == index ? 32'h00000000 : _GEN_776);
	wire [31:0] _GEN_778 = (10'h30a == index ? 32'h00000000 : _GEN_777);
	wire [31:0] _GEN_779 = (10'h30b == index ? 32'h00000000 : _GEN_778);
	wire [31:0] _GEN_780 = (10'h30c == index ? 32'h00000000 : _GEN_779);
	wire [31:0] _GEN_781 = (10'h30d == index ? 32'h00000000 : _GEN_780);
	wire [31:0] _GEN_782 = (10'h30e == index ? 32'h00000000 : _GEN_781);
	wire [31:0] _GEN_783 = (10'h30f == index ? 32'h00000000 : _GEN_782);
	wire [31:0] _GEN_784 = (10'h310 == index ? 32'h00000000 : _GEN_783);
	wire [31:0] _GEN_785 = (10'h311 == index ? 32'h00000000 : _GEN_784);
	wire [31:0] _GEN_786 = (10'h312 == index ? 32'h00000000 : _GEN_785);
	wire [31:0] _GEN_787 = (10'h313 == index ? 32'h00000000 : _GEN_786);
	wire [31:0] _GEN_788 = (10'h314 == index ? 32'h00000000 : _GEN_787);
	wire [31:0] _GEN_789 = (10'h315 == index ? 32'h00000000 : _GEN_788);
	wire [31:0] _GEN_790 = (10'h316 == index ? 32'h00000000 : _GEN_789);
	wire [31:0] _GEN_791 = (10'h317 == index ? 32'h00000000 : _GEN_790);
	wire [31:0] _GEN_792 = (10'h318 == index ? 32'h00000000 : _GEN_791);
	wire [31:0] _GEN_793 = (10'h319 == index ? 32'h00000000 : _GEN_792);
	wire [31:0] _GEN_794 = (10'h31a == index ? 32'h00000000 : _GEN_793);
	wire [31:0] _GEN_795 = (10'h31b == index ? 32'h00000000 : _GEN_794);
	wire [31:0] _GEN_796 = (10'h31c == index ? 32'h00000000 : _GEN_795);
	wire [31:0] _GEN_797 = (10'h31d == index ? 32'h00000000 : _GEN_796);
	wire [31:0] _GEN_798 = (10'h31e == index ? 32'h00000000 : _GEN_797);
	wire [31:0] _GEN_799 = (10'h31f == index ? 32'h00000000 : _GEN_798);
	wire [31:0] _GEN_800 = (10'h320 == index ? 32'h00000000 : _GEN_799);
	wire [31:0] _GEN_801 = (10'h321 == index ? 32'h00000000 : _GEN_800);
	wire [31:0] _GEN_802 = (10'h322 == index ? 32'h00000000 : _GEN_801);
	wire [31:0] _GEN_803 = (10'h323 == index ? 32'h00000000 : _GEN_802);
	wire [31:0] _GEN_804 = (10'h324 == index ? 32'h00000000 : _GEN_803);
	wire [31:0] _GEN_805 = (10'h325 == index ? 32'h00000000 : _GEN_804);
	wire [31:0] _GEN_806 = (10'h326 == index ? 32'h00000000 : _GEN_805);
	wire [31:0] _GEN_807 = (10'h327 == index ? 32'h00000000 : _GEN_806);
	wire [31:0] _GEN_808 = (10'h328 == index ? 32'h00000000 : _GEN_807);
	wire [31:0] _GEN_809 = (10'h329 == index ? 32'h00000000 : _GEN_808);
	wire [31:0] _GEN_810 = (10'h32a == index ? 32'h00000000 : _GEN_809);
	wire [31:0] _GEN_811 = (10'h32b == index ? 32'h00000000 : _GEN_810);
	wire [31:0] _GEN_812 = (10'h32c == index ? 32'h00000000 : _GEN_811);
	wire [31:0] _GEN_813 = (10'h32d == index ? 32'h00000000 : _GEN_812);
	wire [31:0] _GEN_814 = (10'h32e == index ? 32'h00000000 : _GEN_813);
	wire [31:0] _GEN_815 = (10'h32f == index ? 32'h00000000 : _GEN_814);
	wire [31:0] _GEN_816 = (10'h330 == index ? 32'h00000000 : _GEN_815);
	wire [31:0] _GEN_817 = (10'h331 == index ? 32'h00000000 : _GEN_816);
	wire [31:0] _GEN_818 = (10'h332 == index ? 32'h00000000 : _GEN_817);
	wire [31:0] _GEN_819 = (10'h333 == index ? 32'h00000000 : _GEN_818);
	wire [31:0] _GEN_820 = (10'h334 == index ? 32'h00000000 : _GEN_819);
	wire [31:0] _GEN_821 = (10'h335 == index ? 32'h00000000 : _GEN_820);
	wire [31:0] _GEN_822 = (10'h336 == index ? 32'h00000000 : _GEN_821);
	wire [31:0] _GEN_823 = (10'h337 == index ? 32'h00000000 : _GEN_822);
	wire [31:0] _GEN_824 = (10'h338 == index ? 32'h00000000 : _GEN_823);
	wire [31:0] _GEN_825 = (10'h339 == index ? 32'h00000000 : _GEN_824);
	wire [31:0] _GEN_826 = (10'h33a == index ? 32'h00000000 : _GEN_825);
	wire [31:0] _GEN_827 = (10'h33b == index ? 32'h00000000 : _GEN_826);
	wire [31:0] _GEN_828 = (10'h33c == index ? 32'h00000000 : _GEN_827);
	wire [31:0] _GEN_829 = (10'h33d == index ? 32'h00000000 : _GEN_828);
	wire [31:0] _GEN_830 = (10'h33e == index ? 32'h00000000 : _GEN_829);
	wire [31:0] _GEN_831 = (10'h33f == index ? 32'h00000000 : _GEN_830);
	wire [31:0] _GEN_832 = (10'h340 == index ? 32'h00000000 : _GEN_831);
	wire [31:0] _GEN_833 = (10'h341 == index ? 32'h00000000 : _GEN_832);
	wire [31:0] _GEN_834 = (10'h342 == index ? 32'h00000000 : _GEN_833);
	wire [31:0] _GEN_835 = (10'h343 == index ? 32'h00000000 : _GEN_834);
	wire [31:0] _GEN_836 = (10'h344 == index ? 32'h00000000 : _GEN_835);
	wire [31:0] _GEN_837 = (10'h345 == index ? 32'h00000000 : _GEN_836);
	wire [31:0] _GEN_838 = (10'h346 == index ? 32'h00000000 : _GEN_837);
	wire [31:0] _GEN_839 = (10'h347 == index ? 32'h00000000 : _GEN_838);
	wire [31:0] _GEN_840 = (10'h348 == index ? 32'h00000000 : _GEN_839);
	wire [31:0] _GEN_841 = (10'h349 == index ? 32'h00000000 : _GEN_840);
	wire [31:0] _GEN_842 = (10'h34a == index ? 32'h00000000 : _GEN_841);
	wire [31:0] _GEN_843 = (10'h34b == index ? 32'h00000000 : _GEN_842);
	wire [31:0] _GEN_844 = (10'h34c == index ? 32'h00000000 : _GEN_843);
	wire [31:0] _GEN_845 = (10'h34d == index ? 32'h00000000 : _GEN_844);
	wire [31:0] _GEN_846 = (10'h34e == index ? 32'h00000000 : _GEN_845);
	wire [31:0] _GEN_847 = (10'h34f == index ? 32'h00000000 : _GEN_846);
	wire [31:0] _GEN_848 = (10'h350 == index ? 32'h00000000 : _GEN_847);
	wire [31:0] _GEN_849 = (10'h351 == index ? 32'h00000000 : _GEN_848);
	wire [31:0] _GEN_850 = (10'h352 == index ? 32'h00000000 : _GEN_849);
	wire [31:0] _GEN_851 = (10'h353 == index ? 32'h00000000 : _GEN_850);
	wire [31:0] _GEN_852 = (10'h354 == index ? 32'h00000000 : _GEN_851);
	wire [31:0] _GEN_853 = (10'h355 == index ? 32'h00000000 : _GEN_852);
	wire [31:0] _GEN_854 = (10'h356 == index ? 32'h00000000 : _GEN_853);
	wire [31:0] _GEN_855 = (10'h357 == index ? 32'h00000000 : _GEN_854);
	wire [31:0] _GEN_856 = (10'h358 == index ? 32'h00000000 : _GEN_855);
	wire [31:0] _GEN_857 = (10'h359 == index ? 32'h00000000 : _GEN_856);
	wire [31:0] _GEN_858 = (10'h35a == index ? 32'h00000000 : _GEN_857);
	wire [31:0] _GEN_859 = (10'h35b == index ? 32'h00000000 : _GEN_858);
	wire [31:0] _GEN_860 = (10'h35c == index ? 32'h00000000 : _GEN_859);
	wire [31:0] _GEN_861 = (10'h35d == index ? 32'h00000000 : _GEN_860);
	wire [31:0] _GEN_862 = (10'h35e == index ? 32'h00000000 : _GEN_861);
	wire [31:0] _GEN_863 = (10'h35f == index ? 32'h00000000 : _GEN_862);
	wire [31:0] _GEN_864 = (10'h360 == index ? 32'h00000000 : _GEN_863);
	wire [31:0] _GEN_865 = (10'h361 == index ? 32'h00000000 : _GEN_864);
	wire [31:0] _GEN_866 = (10'h362 == index ? 32'h00000000 : _GEN_865);
	wire [31:0] _GEN_867 = (10'h363 == index ? 32'h00000000 : _GEN_866);
	wire [31:0] _GEN_868 = (10'h364 == index ? 32'h00000000 : _GEN_867);
	wire [31:0] _GEN_869 = (10'h365 == index ? 32'h00000000 : _GEN_868);
	wire [31:0] _GEN_870 = (10'h366 == index ? 32'h00000000 : _GEN_869);
	wire [31:0] _GEN_871 = (10'h367 == index ? 32'h00000000 : _GEN_870);
	wire [31:0] _GEN_872 = (10'h368 == index ? 32'h00000000 : _GEN_871);
	wire [31:0] _GEN_873 = (10'h369 == index ? 32'h00000000 : _GEN_872);
	wire [31:0] _GEN_874 = (10'h36a == index ? 32'h00000000 : _GEN_873);
	wire [31:0] _GEN_875 = (10'h36b == index ? 32'h00000000 : _GEN_874);
	wire [31:0] _GEN_876 = (10'h36c == index ? 32'h00000000 : _GEN_875);
	wire [31:0] _GEN_877 = (10'h36d == index ? 32'h00000000 : _GEN_876);
	wire [31:0] _GEN_878 = (10'h36e == index ? 32'h00000000 : _GEN_877);
	wire [31:0] _GEN_879 = (10'h36f == index ? 32'h00000000 : _GEN_878);
	wire [31:0] _GEN_880 = (10'h370 == index ? 32'h00000000 : _GEN_879);
	wire [31:0] _GEN_881 = (10'h371 == index ? 32'h00000000 : _GEN_880);
	wire [31:0] _GEN_882 = (10'h372 == index ? 32'h00000000 : _GEN_881);
	wire [31:0] _GEN_883 = (10'h373 == index ? 32'h00000000 : _GEN_882);
	wire [31:0] _GEN_884 = (10'h374 == index ? 32'h00000000 : _GEN_883);
	wire [31:0] _GEN_885 = (10'h375 == index ? 32'h00000000 : _GEN_884);
	wire [31:0] _GEN_886 = (10'h376 == index ? 32'h00000000 : _GEN_885);
	wire [31:0] _GEN_887 = (10'h377 == index ? 32'h00000000 : _GEN_886);
	wire [31:0] _GEN_888 = (10'h378 == index ? 32'h00000000 : _GEN_887);
	wire [31:0] _GEN_889 = (10'h379 == index ? 32'h00000000 : _GEN_888);
	wire [31:0] _GEN_890 = (10'h37a == index ? 32'h00000000 : _GEN_889);
	wire [31:0] _GEN_891 = (10'h37b == index ? 32'h00000000 : _GEN_890);
	wire [31:0] _GEN_892 = (10'h37c == index ? 32'h00000000 : _GEN_891);
	wire [31:0] _GEN_893 = (10'h37d == index ? 32'h00000000 : _GEN_892);
	wire [31:0] _GEN_894 = (10'h37e == index ? 32'h00000000 : _GEN_893);
	wire [31:0] _GEN_895 = (10'h37f == index ? 32'h00000000 : _GEN_894);
	wire [31:0] _GEN_896 = (10'h380 == index ? 32'h00000000 : _GEN_895);
	wire [31:0] _GEN_897 = (10'h381 == index ? 32'h00000000 : _GEN_896);
	wire [31:0] _GEN_898 = (10'h382 == index ? 32'h00000000 : _GEN_897);
	wire [31:0] _GEN_899 = (10'h383 == index ? 32'h00000000 : _GEN_898);
	wire [31:0] _GEN_900 = (10'h384 == index ? 32'h00000000 : _GEN_899);
	wire [31:0] _GEN_901 = (10'h385 == index ? 32'h00000000 : _GEN_900);
	wire [31:0] _GEN_902 = (10'h386 == index ? 32'h00000000 : _GEN_901);
	wire [31:0] _GEN_903 = (10'h387 == index ? 32'h00000000 : _GEN_902);
	wire [31:0] _GEN_904 = (10'h388 == index ? 32'h00000000 : _GEN_903);
	wire [31:0] _GEN_905 = (10'h389 == index ? 32'h00000000 : _GEN_904);
	wire [31:0] _GEN_906 = (10'h38a == index ? 32'h00000000 : _GEN_905);
	wire [31:0] _GEN_907 = (10'h38b == index ? 32'h00000000 : _GEN_906);
	wire [31:0] _GEN_908 = (10'h38c == index ? 32'h00000000 : _GEN_907);
	wire [31:0] _GEN_909 = (10'h38d == index ? 32'h00000000 : _GEN_908);
	wire [31:0] _GEN_910 = (10'h38e == index ? 32'h00000000 : _GEN_909);
	wire [31:0] _GEN_911 = (10'h38f == index ? 32'h00000000 : _GEN_910);
	wire [31:0] _GEN_912 = (10'h390 == index ? 32'h00000000 : _GEN_911);
	wire [31:0] _GEN_913 = (10'h391 == index ? 32'h00000000 : _GEN_912);
	wire [31:0] _GEN_914 = (10'h392 == index ? 32'h00000000 : _GEN_913);
	wire [31:0] _GEN_915 = (10'h393 == index ? 32'h00000000 : _GEN_914);
	wire [31:0] _GEN_916 = (10'h394 == index ? 32'h00000000 : _GEN_915);
	wire [31:0] _GEN_917 = (10'h395 == index ? 32'h00000000 : _GEN_916);
	wire [31:0] _GEN_918 = (10'h396 == index ? 32'h00000000 : _GEN_917);
	wire [31:0] _GEN_919 = (10'h397 == index ? 32'h00000000 : _GEN_918);
	wire [31:0] _GEN_920 = (10'h398 == index ? 32'h00000000 : _GEN_919);
	wire [31:0] _GEN_921 = (10'h399 == index ? 32'h00000000 : _GEN_920);
	wire [31:0] _GEN_922 = (10'h39a == index ? 32'h00000000 : _GEN_921);
	wire [31:0] _GEN_923 = (10'h39b == index ? 32'h00000000 : _GEN_922);
	wire [31:0] _GEN_924 = (10'h39c == index ? 32'h00000000 : _GEN_923);
	wire [31:0] _GEN_925 = (10'h39d == index ? 32'h00000000 : _GEN_924);
	wire [31:0] _GEN_926 = (10'h39e == index ? 32'h00000000 : _GEN_925);
	wire [31:0] _GEN_927 = (10'h39f == index ? 32'h00000000 : _GEN_926);
	wire [31:0] _GEN_928 = (10'h3a0 == index ? 32'h00000000 : _GEN_927);
	wire [31:0] _GEN_929 = (10'h3a1 == index ? 32'h00000000 : _GEN_928);
	wire [31:0] _GEN_930 = (10'h3a2 == index ? 32'h00000000 : _GEN_929);
	wire [31:0] _GEN_931 = (10'h3a3 == index ? 32'h00000000 : _GEN_930);
	wire [31:0] _GEN_932 = (10'h3a4 == index ? 32'h00000000 : _GEN_931);
	wire [31:0] _GEN_933 = (10'h3a5 == index ? 32'h00000000 : _GEN_932);
	wire [31:0] _GEN_934 = (10'h3a6 == index ? 32'h00000000 : _GEN_933);
	wire [31:0] _GEN_935 = (10'h3a7 == index ? 32'h00000000 : _GEN_934);
	wire [31:0] _GEN_936 = (10'h3a8 == index ? 32'h00000000 : _GEN_935);
	wire [31:0] _GEN_937 = (10'h3a9 == index ? 32'h00000000 : _GEN_936);
	wire [31:0] _GEN_938 = (10'h3aa == index ? 32'h00000000 : _GEN_937);
	wire [31:0] _GEN_939 = (10'h3ab == index ? 32'h00000000 : _GEN_938);
	wire [31:0] _GEN_940 = (10'h3ac == index ? 32'h00000000 : _GEN_939);
	wire [31:0] _GEN_941 = (10'h3ad == index ? 32'h00000000 : _GEN_940);
	wire [31:0] _GEN_942 = (10'h3ae == index ? 32'h00000000 : _GEN_941);
	wire [31:0] _GEN_943 = (10'h3af == index ? 32'h00000000 : _GEN_942);
	wire [31:0] _GEN_944 = (10'h3b0 == index ? 32'h00000000 : _GEN_943);
	wire [31:0] _GEN_945 = (10'h3b1 == index ? 32'h00000000 : _GEN_944);
	wire [31:0] _GEN_946 = (10'h3b2 == index ? 32'h00000000 : _GEN_945);
	wire [31:0] _GEN_947 = (10'h3b3 == index ? 32'h00000000 : _GEN_946);
	wire [31:0] _GEN_948 = (10'h3b4 == index ? 32'h00000000 : _GEN_947);
	wire [31:0] _GEN_949 = (10'h3b5 == index ? 32'h00000000 : _GEN_948);
	wire [31:0] _GEN_950 = (10'h3b6 == index ? 32'h00000000 : _GEN_949);
	wire [31:0] _GEN_951 = (10'h3b7 == index ? 32'h00000000 : _GEN_950);
	wire [31:0] _GEN_952 = (10'h3b8 == index ? 32'h00000000 : _GEN_951);
	wire [31:0] _GEN_953 = (10'h3b9 == index ? 32'h00000000 : _GEN_952);
	wire [31:0] _GEN_954 = (10'h3ba == index ? 32'h00000000 : _GEN_953);
	wire [31:0] _GEN_955 = (10'h3bb == index ? 32'h00000000 : _GEN_954);
	wire [31:0] _GEN_956 = (10'h3bc == index ? 32'h00000000 : _GEN_955);
	wire [31:0] _GEN_957 = (10'h3bd == index ? 32'h00000000 : _GEN_956);
	wire [31:0] _GEN_958 = (10'h3be == index ? 32'h00000000 : _GEN_957);
	wire [31:0] _GEN_959 = (10'h3bf == index ? 32'h00000000 : _GEN_958);
	wire [31:0] _GEN_960 = (10'h3c0 == index ? 32'h00000000 : _GEN_959);
	wire [31:0] _GEN_961 = (10'h3c1 == index ? 32'h00000000 : _GEN_960);
	wire [31:0] _GEN_962 = (10'h3c2 == index ? 32'h00000000 : _GEN_961);
	wire [31:0] _GEN_963 = (10'h3c3 == index ? 32'h00000000 : _GEN_962);
	wire [31:0] _GEN_964 = (10'h3c4 == index ? 32'h00000000 : _GEN_963);
	wire [31:0] _GEN_965 = (10'h3c5 == index ? 32'h00000000 : _GEN_964);
	wire [31:0] _GEN_966 = (10'h3c6 == index ? 32'h00000000 : _GEN_965);
	wire [31:0] _GEN_967 = (10'h3c7 == index ? 32'h00000000 : _GEN_966);
	wire [31:0] _GEN_968 = (10'h3c8 == index ? 32'h00000000 : _GEN_967);
	wire [31:0] _GEN_969 = (10'h3c9 == index ? 32'h00000000 : _GEN_968);
	wire [31:0] _GEN_970 = (10'h3ca == index ? 32'h00000000 : _GEN_969);
	wire [31:0] _GEN_971 = (10'h3cb == index ? 32'h00000000 : _GEN_970);
	wire [31:0] _GEN_972 = (10'h3cc == index ? 32'h00000000 : _GEN_971);
	wire [31:0] _GEN_973 = (10'h3cd == index ? 32'h00000000 : _GEN_972);
	wire [31:0] _GEN_974 = (10'h3ce == index ? 32'h00000000 : _GEN_973);
	wire [31:0] _GEN_975 = (10'h3cf == index ? 32'h00000000 : _GEN_974);
	wire [31:0] _GEN_976 = (10'h3d0 == index ? 32'h00000000 : _GEN_975);
	wire [31:0] _GEN_977 = (10'h3d1 == index ? 32'h00000000 : _GEN_976);
	wire [31:0] _GEN_978 = (10'h3d2 == index ? 32'h00000000 : _GEN_977);
	wire [31:0] _GEN_979 = (10'h3d3 == index ? 32'h00000000 : _GEN_978);
	wire [31:0] _GEN_980 = (10'h3d4 == index ? 32'h00000000 : _GEN_979);
	wire [31:0] _GEN_981 = (10'h3d5 == index ? 32'h00000000 : _GEN_980);
	wire [31:0] _GEN_982 = (10'h3d6 == index ? 32'h00000000 : _GEN_981);
	wire [31:0] _GEN_983 = (10'h3d7 == index ? 32'h00000000 : _GEN_982);
	wire [31:0] _GEN_984 = (10'h3d8 == index ? 32'h00000000 : _GEN_983);
	wire [31:0] _GEN_985 = (10'h3d9 == index ? 32'h00000000 : _GEN_984);
	wire [31:0] _GEN_986 = (10'h3da == index ? 32'h00000000 : _GEN_985);
	wire [31:0] _GEN_987 = (10'h3db == index ? 32'h00000000 : _GEN_986);
	wire [31:0] _GEN_988 = (10'h3dc == index ? 32'h00000000 : _GEN_987);
	wire [31:0] _GEN_989 = (10'h3dd == index ? 32'h00000000 : _GEN_988);
	wire [31:0] _GEN_990 = (10'h3de == index ? 32'h00000000 : _GEN_989);
	wire [31:0] _GEN_991 = (10'h3df == index ? 32'h00000000 : _GEN_990);
	wire [31:0] _GEN_992 = (10'h3e0 == index ? 32'h00000000 : _GEN_991);
	wire [31:0] _GEN_993 = (10'h3e1 == index ? 32'h00000000 : _GEN_992);
	wire [31:0] _GEN_994 = (10'h3e2 == index ? 32'h00000000 : _GEN_993);
	wire [31:0] _GEN_995 = (10'h3e3 == index ? 32'h00000000 : _GEN_994);
	wire [31:0] _GEN_996 = (10'h3e4 == index ? 32'h00000000 : _GEN_995);
	wire [31:0] _GEN_997 = (10'h3e5 == index ? 32'h00000000 : _GEN_996);
	wire [31:0] _GEN_998 = (10'h3e6 == index ? 32'h00000000 : _GEN_997);
	wire [31:0] _GEN_999 = (10'h3e7 == index ? 32'h00000000 : _GEN_998);
	wire [31:0] _GEN_1000 = (10'h3e8 == index ? 32'h00000000 : _GEN_999);
	wire [31:0] _GEN_1001 = (10'h3e9 == index ? 32'h00000000 : _GEN_1000);
	wire [31:0] _GEN_1002 = (10'h3ea == index ? 32'h00000000 : _GEN_1001);
	wire [31:0] _GEN_1003 = (10'h3eb == index ? 32'h00000000 : _GEN_1002);
	wire [31:0] _GEN_1004 = (10'h3ec == index ? 32'h00000000 : _GEN_1003);
	wire [31:0] _GEN_1005 = (10'h3ed == index ? 32'h00000000 : _GEN_1004);
	wire [31:0] _GEN_1006 = (10'h3ee == index ? 32'h00000000 : _GEN_1005);
	wire [31:0] _GEN_1007 = (10'h3ef == index ? 32'h00000000 : _GEN_1006);
	wire [31:0] _GEN_1008 = (10'h3f0 == index ? 32'h00000000 : _GEN_1007);
	wire [31:0] _GEN_1009 = (10'h3f1 == index ? 32'h00000000 : _GEN_1008);
	wire [31:0] _GEN_1010 = (10'h3f2 == index ? 32'h00000000 : _GEN_1009);
	wire [31:0] _GEN_1011 = (10'h3f3 == index ? 32'h00000000 : _GEN_1010);
	wire [31:0] _GEN_1012 = (10'h3f4 == index ? 32'h00000000 : _GEN_1011);
	wire [31:0] _GEN_1013 = (10'h3f5 == index ? 32'h00000000 : _GEN_1012);
	wire [31:0] _GEN_1014 = (10'h3f6 == index ? 32'h00000000 : _GEN_1013);
	wire [31:0] _GEN_1015 = (10'h3f7 == index ? 32'h00000000 : _GEN_1014);
	wire [31:0] _GEN_1016 = (10'h3f8 == index ? 32'h00000000 : _GEN_1015);
	wire [31:0] _GEN_1017 = (10'h3f9 == index ? 32'h00000000 : _GEN_1016);
	wire [31:0] _GEN_1018 = (10'h3fa == index ? 32'h00000000 : _GEN_1017);
	wire [31:0] _GEN_1019 = (10'h3fb == index ? 32'h00000000 : _GEN_1018);
	wire [31:0] _GEN_1020 = (10'h3fc == index ? 32'h00000000 : _GEN_1019);
	wire [31:0] _GEN_1021 = (10'h3fd == index ? 32'h00000000 : _GEN_1020);
	wire [31:0] _GEN_1022 = (10'h3fe == index ? 32'h00000000 : _GEN_1021);
	wire [31:0] _GEN_1023 = (10'h3ff == index ? 32'h00000000 : _GEN_1022);
	TLMonitor_43 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	assign auto_in_a_ready = auto_in_d_ready;
	assign auto_in_d_valid = auto_in_a_valid;
	assign auto_in_d_bits_size = auto_in_a_bits_size;
	assign auto_in_d_bits_source = auto_in_a_bits_source;
	assign auto_in_d_bits_data = (|high ? 32'h00000000 : _GEN_1023);
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_in_d_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = auto_in_a_valid;
	assign monitor_io_in_d_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_d_bits_source = auto_in_a_bits_source;
endmodule
module ClockSinkDomain_1 (
	auto_bootrom_in_a_ready,
	auto_bootrom_in_a_valid,
	auto_bootrom_in_a_bits_opcode,
	auto_bootrom_in_a_bits_param,
	auto_bootrom_in_a_bits_size,
	auto_bootrom_in_a_bits_source,
	auto_bootrom_in_a_bits_address,
	auto_bootrom_in_a_bits_mask,
	auto_bootrom_in_a_bits_corrupt,
	auto_bootrom_in_d_ready,
	auto_bootrom_in_d_valid,
	auto_bootrom_in_d_bits_size,
	auto_bootrom_in_d_bits_source,
	auto_bootrom_in_d_bits_data,
	auto_clock_in_clock,
	auto_clock_in_reset
);
	output wire auto_bootrom_in_a_ready;
	input auto_bootrom_in_a_valid;
	input [2:0] auto_bootrom_in_a_bits_opcode;
	input [2:0] auto_bootrom_in_a_bits_param;
	input [1:0] auto_bootrom_in_a_bits_size;
	input [7:0] auto_bootrom_in_a_bits_source;
	input [16:0] auto_bootrom_in_a_bits_address;
	input [3:0] auto_bootrom_in_a_bits_mask;
	input auto_bootrom_in_a_bits_corrupt;
	input auto_bootrom_in_d_ready;
	output wire auto_bootrom_in_d_valid;
	output wire [1:0] auto_bootrom_in_d_bits_size;
	output wire [7:0] auto_bootrom_in_d_bits_source;
	output wire [31:0] auto_bootrom_in_d_bits_data;
	input auto_clock_in_clock;
	input auto_clock_in_reset;
	wire bootrom_clock;
	wire bootrom_reset;
	wire bootrom_auto_in_a_ready;
	wire bootrom_auto_in_a_valid;
	wire [2:0] bootrom_auto_in_a_bits_opcode;
	wire [2:0] bootrom_auto_in_a_bits_param;
	wire [1:0] bootrom_auto_in_a_bits_size;
	wire [7:0] bootrom_auto_in_a_bits_source;
	wire [16:0] bootrom_auto_in_a_bits_address;
	wire [3:0] bootrom_auto_in_a_bits_mask;
	wire bootrom_auto_in_a_bits_corrupt;
	wire bootrom_auto_in_d_ready;
	wire bootrom_auto_in_d_valid;
	wire [1:0] bootrom_auto_in_d_bits_size;
	wire [7:0] bootrom_auto_in_d_bits_source;
	wire [31:0] bootrom_auto_in_d_bits_data;
	TLROM bootrom(
		.clock(bootrom_clock),
		.reset(bootrom_reset),
		.auto_in_a_ready(bootrom_auto_in_a_ready),
		.auto_in_a_valid(bootrom_auto_in_a_valid),
		.auto_in_a_bits_opcode(bootrom_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(bootrom_auto_in_a_bits_param),
		.auto_in_a_bits_size(bootrom_auto_in_a_bits_size),
		.auto_in_a_bits_source(bootrom_auto_in_a_bits_source),
		.auto_in_a_bits_address(bootrom_auto_in_a_bits_address),
		.auto_in_a_bits_mask(bootrom_auto_in_a_bits_mask),
		.auto_in_a_bits_corrupt(bootrom_auto_in_a_bits_corrupt),
		.auto_in_d_ready(bootrom_auto_in_d_ready),
		.auto_in_d_valid(bootrom_auto_in_d_valid),
		.auto_in_d_bits_size(bootrom_auto_in_d_bits_size),
		.auto_in_d_bits_source(bootrom_auto_in_d_bits_source),
		.auto_in_d_bits_data(bootrom_auto_in_d_bits_data)
	);
	assign auto_bootrom_in_a_ready = bootrom_auto_in_a_ready;
	assign auto_bootrom_in_d_valid = bootrom_auto_in_d_valid;
	assign auto_bootrom_in_d_bits_size = bootrom_auto_in_d_bits_size;
	assign auto_bootrom_in_d_bits_source = bootrom_auto_in_d_bits_source;
	assign auto_bootrom_in_d_bits_data = bootrom_auto_in_d_bits_data;
	assign bootrom_clock = auto_clock_in_clock;
	assign bootrom_reset = auto_clock_in_reset;
	assign bootrom_auto_in_a_valid = auto_bootrom_in_a_valid;
	assign bootrom_auto_in_a_bits_opcode = auto_bootrom_in_a_bits_opcode;
	assign bootrom_auto_in_a_bits_param = auto_bootrom_in_a_bits_param;
	assign bootrom_auto_in_a_bits_size = auto_bootrom_in_a_bits_size;
	assign bootrom_auto_in_a_bits_source = auto_bootrom_in_a_bits_source;
	assign bootrom_auto_in_a_bits_address = auto_bootrom_in_a_bits_address;
	assign bootrom_auto_in_a_bits_mask = auto_bootrom_in_a_bits_mask;
	assign bootrom_auto_in_a_bits_corrupt = auto_bootrom_in_a_bits_corrupt;
	assign bootrom_auto_in_d_ready = auto_bootrom_in_d_ready;
endmodule
module TLMonitor_44 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [28:0] io_in_a_bits_address;
	input [7:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [28:0] _GEN_71 = {23'd0, is_aligned_mask};
	wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 29'h00000000;
	wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0];
	wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount;
	wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h3;
	wire mask_size = mask_sizeOH[2];
	wire mask_bit = io_in_a_bits_address[2];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[1];
	wire mask_bit_1 = io_in_a_bits_address[1];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire mask_size_2 = mask_sizeOH[0];
	wire mask_bit_2 = io_in_a_bits_address[0];
	wire mask_nbit_2 = ~mask_bit_2;
	wire mask_eq_6 = mask_eq_2 & mask_nbit_2;
	wire mask_acc_6 = mask_acc_2 | (mask_size_2 & mask_eq_6);
	wire mask_eq_7 = mask_eq_2 & mask_bit_2;
	wire mask_acc_7 = mask_acc_2 | (mask_size_2 & mask_eq_7);
	wire mask_eq_8 = mask_eq_3 & mask_nbit_2;
	wire mask_acc_8 = mask_acc_3 | (mask_size_2 & mask_eq_8);
	wire mask_eq_9 = mask_eq_3 & mask_bit_2;
	wire mask_acc_9 = mask_acc_3 | (mask_size_2 & mask_eq_9);
	wire mask_eq_10 = mask_eq_4 & mask_nbit_2;
	wire mask_acc_10 = mask_acc_4 | (mask_size_2 & mask_eq_10);
	wire mask_eq_11 = mask_eq_4 & mask_bit_2;
	wire mask_acc_11 = mask_acc_4 | (mask_size_2 & mask_eq_11);
	wire mask_eq_12 = mask_eq_5 & mask_nbit_2;
	wire mask_acc_12 = mask_acc_5 | (mask_size_2 & mask_eq_12);
	wire mask_eq_13 = mask_eq_5 & mask_bit_2;
	wire mask_acc_13 = mask_acc_5 | (mask_size_2 & mask_eq_13);
	wire [7:0] mask = {mask_acc_13, mask_acc_12, mask_acc_11, mask_acc_10, mask_acc_9, mask_acc_8, mask_acc_7, mask_acc_6};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [28:0] _T_56 = io_in_a_bits_address ^ 29'h00020000;
	wire [29:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [29:0] _T_59 = $signed(_T_57) & -30'sh00010000;
	wire _T_60 = $signed(_T_59) == 30'sh00000000;
	wire [28:0] _T_61 = io_in_a_bits_address ^ 29'h10000000;
	wire [29:0] _T_62 = {1'b0, $signed(_T_61)};
	wire [29:0] _T_64 = $signed(_T_62) & -30'sh00001000;
	wire _T_65 = $signed(_T_64) == 30'sh00000000;
	wire _T_66 = _T_60 | _T_65;
	wire _T_104 = io_in_a_bits_param <= 3'h2;
	wire [7:0] _T_108 = ~io_in_a_bits_mask;
	wire _T_109 = _T_108 == 8'h00;
	wire _T_113 = ~io_in_a_bits_corrupt;
	wire _T_117 = io_in_a_bits_opcode == 3'h7;
	wire _T_183 = io_in_a_bits_param != 3'h0;
	wire _T_196 = io_in_a_bits_opcode == 3'h4;
	wire _T_213 = io_in_a_bits_size <= 3'h6;
	wire _T_227 = _T_213 & _T_66;
	wire _T_238 = io_in_a_bits_param == 3'h0;
	wire _T_242 = io_in_a_bits_mask == mask;
	wire _T_250 = io_in_a_bits_opcode == 3'h0;
	wire _T_272 = _T_213 & _T_65;
	wire _T_282 = source_ok & _T_272;
	wire _T_300 = io_in_a_bits_opcode == 3'h1;
	wire [7:0] _T_346 = ~mask;
	wire [7:0] _T_347 = io_in_a_bits_mask & _T_346;
	wire _T_348 = _T_347 == 8'h00;
	wire _T_352 = io_in_a_bits_opcode == 3'h2;
	wire _T_389 = io_in_a_bits_param <= 3'h4;
	wire _T_397 = io_in_a_bits_opcode == 3'h3;
	wire _T_434 = io_in_a_bits_param <= 3'h3;
	wire _T_442 = io_in_a_bits_opcode == 3'h5;
	wire _T_479 = io_in_a_bits_param <= 3'h1;
	wire _T_491 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_495 = io_in_d_bits_opcode == 3'h6;
	wire _T_499 = io_in_d_bits_size >= 3'h3;
	wire _T_503 = io_in_d_bits_param == 2'h0;
	wire _T_507 = ~io_in_d_bits_corrupt;
	wire _T_511 = ~io_in_d_bits_denied;
	wire _T_515 = io_in_d_bits_opcode == 3'h4;
	wire _T_526 = io_in_d_bits_param <= 2'h2;
	wire _T_530 = io_in_d_bits_param != 2'h2;
	wire _T_543 = io_in_d_bits_opcode == 3'h5;
	wire _T_563 = _T_511 | io_in_d_bits_corrupt;
	wire _T_572 = io_in_d_bits_opcode == 3'h0;
	wire _T_589 = io_in_d_bits_opcode == 3'h1;
	wire _T_607 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [2:0] a_first_counter;
	wire [2:0] a_first_counter1 = a_first_counter - 3'h1;
	wire a_first = a_first_counter == 3'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [28:0] address;
	wire _T_637 = io_in_a_valid & ~a_first;
	wire _T_638 = io_in_a_bits_opcode == opcode;
	wire _T_642 = io_in_a_bits_param == param;
	wire _T_646 = io_in_a_bits_size == size;
	wire _T_650 = io_in_a_bits_source == source;
	wire _T_654 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [2:0] d_first_counter;
	wire [2:0] d_first_counter1 = d_first_counter - 3'h1;
	wire d_first = d_first_counter == 3'h0;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_661 = io_in_d_valid & ~d_first;
	wire _T_662 = io_in_d_bits_opcode == opcode_1;
	wire _T_666 = io_in_d_bits_param == param_1;
	wire _T_670 = io_in_d_bits_size == size_1;
	wire _T_674 = io_in_d_bits_source == source_1;
	wire _T_678 = io_in_d_bits_sink == sink;
	wire _T_682 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [2:0] a_first_counter_1;
	wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1;
	wire a_first_1 = a_first_counter_1 == 3'h0;
	reg [2:0] d_first_counter_1;
	wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1;
	wire d_first_1 = d_first_counter_1 == 3'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_688 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire _T_691 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_693 = inflight >> io_in_a_bits_source;
	wire _T_695 = ~_T_693[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_699 = io_in_d_valid & d_first_1;
	wire _T_701 = ~_T_495;
	wire _T_702 = (io_in_d_valid & d_first_1) & ~_T_495;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_701 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_701 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_688 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_712 = inflight >> io_in_d_bits_source;
	wire _T_714 = _T_712[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_719 = io_in_d_bits_opcode == _GEN_40;
	wire _T_720 = (io_in_d_bits_opcode == _GEN_32) | _T_719;
	wire _T_724 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_731 = io_in_d_bits_opcode == _GEN_56;
	wire _T_732 = (io_in_d_bits_opcode == _GEN_48) | _T_731;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_736 = _GEN_82 == a_size_lookup;
	wire _T_746 = (((_T_699 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_701;
	wire _T_748 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_757 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [2:0] d_first_counter_2;
	wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1;
	wire d_first_2 = d_first_counter_2 == 3'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_783 = (io_in_d_valid & d_first_2) & _T_495;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_495 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_495 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_791 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_801 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_821 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 3'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 3'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 3'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 3'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 3'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 3'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 3'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 3'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 3'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 3'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module HellaPeekingArbiter (
	clock,
	reset,
	io_in_1_ready,
	io_in_1_valid,
	io_in_1_bits_opcode,
	io_in_1_bits_param,
	io_in_1_bits_size,
	io_in_1_bits_source,
	io_in_1_bits_data,
	io_in_1_bits_corrupt,
	io_in_1_bits_union,
	io_in_1_bits_last,
	io_in_4_ready,
	io_in_4_valid,
	io_in_4_bits_opcode,
	io_in_4_bits_param,
	io_in_4_bits_size,
	io_in_4_bits_source,
	io_in_4_bits_address,
	io_in_4_bits_data,
	io_in_4_bits_corrupt,
	io_in_4_bits_union,
	io_in_4_bits_last,
	io_out_ready,
	io_out_valid,
	io_out_bits_chanId,
	io_out_bits_opcode,
	io_out_bits_param,
	io_out_bits_size,
	io_out_bits_source,
	io_out_bits_address,
	io_out_bits_data,
	io_out_bits_corrupt,
	io_out_bits_union,
	io_out_bits_last
);
	input clock;
	input reset;
	output wire io_in_1_ready;
	input io_in_1_valid;
	input [2:0] io_in_1_bits_opcode;
	input [2:0] io_in_1_bits_param;
	input [3:0] io_in_1_bits_size;
	input [2:0] io_in_1_bits_source;
	input [63:0] io_in_1_bits_data;
	input io_in_1_bits_corrupt;
	input [7:0] io_in_1_bits_union;
	input io_in_1_bits_last;
	output wire io_in_4_ready;
	input io_in_4_valid;
	input [2:0] io_in_4_bits_opcode;
	input [2:0] io_in_4_bits_param;
	input [3:0] io_in_4_bits_size;
	input [2:0] io_in_4_bits_source;
	input [31:0] io_in_4_bits_address;
	input [63:0] io_in_4_bits_data;
	input io_in_4_bits_corrupt;
	input [7:0] io_in_4_bits_union;
	input io_in_4_bits_last;
	input io_out_ready;
	output wire io_out_valid;
	output wire [2:0] io_out_bits_chanId;
	output wire [2:0] io_out_bits_opcode;
	output wire [2:0] io_out_bits_param;
	output wire [3:0] io_out_bits_size;
	output wire [2:0] io_out_bits_source;
	output wire [31:0] io_out_bits_address;
	output wire [63:0] io_out_bits_data;
	output wire io_out_bits_corrupt;
	output wire [7:0] io_out_bits_union;
	output wire io_out_bits_last;
	reg [2:0] lockIdx;
	reg locked;
	wire [2:0] choice = (io_in_1_valid ? 3'h1 : 3'h4);
	wire [2:0] chosen = (locked ? lockIdx : choice);
	wire _GEN_60 = 3'h1 == chosen;
	wire _GEN_2 = (3'h2 == chosen ? 1'h0 : (3'h1 == chosen) & io_in_1_valid);
	wire _GEN_3 = (3'h3 == chosen ? 1'h0 : _GEN_2);
	wire [2:0] _GEN_6 = (3'h1 == chosen ? 3'h3 : 3'h4);
	wire [2:0] _GEN_7 = (3'h2 == chosen ? 3'h2 : _GEN_6);
	wire [2:0] _GEN_8 = (3'h3 == chosen ? 3'h1 : _GEN_7);
	wire [2:0] _GEN_11 = (3'h1 == chosen ? io_in_1_bits_opcode : 3'h0);
	wire [2:0] _GEN_12 = (3'h2 == chosen ? 3'h0 : _GEN_11);
	wire [2:0] _GEN_13 = (3'h3 == chosen ? 3'h0 : _GEN_12);
	wire [2:0] _GEN_16 = (3'h1 == chosen ? io_in_1_bits_param : 3'h0);
	wire [2:0] _GEN_17 = (3'h2 == chosen ? 3'h0 : _GEN_16);
	wire [2:0] _GEN_18 = (3'h3 == chosen ? 3'h0 : _GEN_17);
	wire [3:0] _GEN_21 = (3'h1 == chosen ? io_in_1_bits_size : 4'h0);
	wire [3:0] _GEN_22 = (3'h2 == chosen ? 4'h0 : _GEN_21);
	wire [3:0] _GEN_23 = (3'h3 == chosen ? 4'h0 : _GEN_22);
	wire [2:0] _GEN_26 = (3'h1 == chosen ? io_in_1_bits_source : 3'h0);
	wire [2:0] _GEN_27 = (3'h2 == chosen ? 3'h0 : _GEN_26);
	wire [2:0] _GEN_28 = (3'h3 == chosen ? 3'h0 : _GEN_27);
	wire [63:0] _GEN_36 = (3'h1 == chosen ? io_in_1_bits_data : 64'h0000000000000000);
	wire [63:0] _GEN_37 = (3'h2 == chosen ? 64'h0000000000000000 : _GEN_36);
	wire [63:0] _GEN_38 = (3'h3 == chosen ? 64'h0000000000000000 : _GEN_37);
	wire _GEN_42 = (3'h2 == chosen ? 1'h0 : _GEN_60 & io_in_1_bits_corrupt);
	wire _GEN_43 = (3'h3 == chosen ? 1'h0 : _GEN_42);
	wire [7:0] _GEN_46 = (3'h1 == chosen ? io_in_1_bits_union : 8'h00);
	wire [7:0] _GEN_47 = (3'h2 == chosen ? 8'h00 : _GEN_46);
	wire [7:0] _GEN_48 = (3'h3 == chosen ? 8'h00 : _GEN_47);
	wire _GEN_51 = (3'h1 == chosen ? io_in_1_bits_last : 1'h1);
	wire _T = io_out_ready & io_out_valid;
	wire _GEN_56 = ~locked | locked;
	assign io_in_1_ready = io_out_ready & (chosen == 3'h1);
	assign io_in_4_ready = io_out_ready & (chosen == 3'h4);
	assign io_out_valid = (3'h4 == chosen ? io_in_4_valid : _GEN_3);
	assign io_out_bits_chanId = (3'h4 == chosen ? 3'h0 : _GEN_8);
	assign io_out_bits_opcode = (3'h4 == chosen ? io_in_4_bits_opcode : _GEN_13);
	assign io_out_bits_param = (3'h4 == chosen ? io_in_4_bits_param : _GEN_18);
	assign io_out_bits_size = (3'h4 == chosen ? io_in_4_bits_size : _GEN_23);
	assign io_out_bits_source = (3'h4 == chosen ? io_in_4_bits_source : _GEN_28);
	assign io_out_bits_address = (3'h4 == chosen ? io_in_4_bits_address : 32'h00000000);
	assign io_out_bits_data = (3'h4 == chosen ? io_in_4_bits_data : _GEN_38);
	assign io_out_bits_corrupt = (3'h4 == chosen ? io_in_4_bits_corrupt : _GEN_43);
	assign io_out_bits_union = (3'h4 == chosen ? io_in_4_bits_union : _GEN_48);
	assign io_out_bits_last = (3'h4 == chosen ? io_in_4_bits_last : (3'h3 == chosen) | ((3'h2 == chosen) | _GEN_51));
	always @(posedge clock) begin
		if (reset)
			lockIdx <= 3'h0;
		else if (_T)
			if (~locked)
				if (io_in_1_valid)
					lockIdx <= 3'h1;
				else
					lockIdx <= 3'h4;
		if (reset)
			locked <= 1'h0;
		else if (_T)
			if (io_out_bits_last)
				locked <= 1'h0;
			else
				locked <= _GEN_56;
	end
endmodule
module GenericSerializer (
	clock,
	reset,
	io_in_ready,
	io_in_valid,
	io_in_bits_chanId,
	io_in_bits_opcode,
	io_in_bits_param,
	io_in_bits_size,
	io_in_bits_source,
	io_in_bits_address,
	io_in_bits_data,
	io_in_bits_corrupt,
	io_in_bits_union,
	io_in_bits_last,
	io_out_ready,
	io_out_valid,
	io_out_bits
);
	input clock;
	input reset;
	output wire io_in_ready;
	input io_in_valid;
	input [2:0] io_in_bits_chanId;
	input [2:0] io_in_bits_opcode;
	input [2:0] io_in_bits_param;
	input [3:0] io_in_bits_size;
	input [2:0] io_in_bits_source;
	input [31:0] io_in_bits_address;
	input [63:0] io_in_bits_data;
	input io_in_bits_corrupt;
	input [7:0] io_in_bits_union;
	input io_in_bits_last;
	input io_out_ready;
	output wire io_out_valid;
	output wire [31:0] io_out_bits;
	reg [121:0] data;
	reg sending;
	wire _T = io_out_ready & io_out_valid;
	reg [1:0] sendCount;
	wire wrap_wrap = sendCount == 2'h3;
	wire [1:0] _wrap_value_T_1 = sendCount + 2'h1;
	wire sendDone = _T & wrap_wrap;
	wire _T_1 = io_in_ready & io_in_valid;
	wire [121:0] _data_T = {io_in_bits_chanId, io_in_bits_opcode, io_in_bits_param, io_in_bits_size, io_in_bits_source, io_in_bits_address, io_in_bits_data, io_in_bits_corrupt, io_in_bits_union, io_in_bits_last};
	wire _GEN_3 = _T_1 | sending;
	wire [121:0] _data_T_1 = {32'd0, data[121:32]};
	assign io_in_ready = ~sending;
	assign io_out_valid = sending;
	assign io_out_bits = data[31:0];
	always @(posedge clock) begin
		if (_T)
			data <= _data_T_1;
		else if (_T_1)
			data <= _data_T;
		if (reset)
			sending <= 1'h0;
		else if (sendDone)
			sending <= 1'h0;
		else
			sending <= _GEN_3;
		if (reset)
			sendCount <= 2'h0;
		else if (_T)
			sendCount <= _wrap_value_T_1;
	end
endmodule
module GenericDeserializer (
	clock,
	reset,
	io_in_ready,
	io_in_valid,
	io_in_bits,
	io_out_ready,
	io_out_valid,
	io_out_bits_chanId,
	io_out_bits_opcode,
	io_out_bits_param,
	io_out_bits_size,
	io_out_bits_source,
	io_out_bits_address,
	io_out_bits_data,
	io_out_bits_corrupt,
	io_out_bits_union
);
	input clock;
	input reset;
	output wire io_in_ready;
	input io_in_valid;
	input [31:0] io_in_bits;
	input io_out_ready;
	output wire io_out_valid;
	output wire [2:0] io_out_bits_chanId;
	output wire [2:0] io_out_bits_opcode;
	output wire [2:0] io_out_bits_param;
	output wire [3:0] io_out_bits_size;
	output wire [2:0] io_out_bits_source;
	output wire [31:0] io_out_bits_address;
	output wire [63:0] io_out_bits_data;
	output wire io_out_bits_corrupt;
	output wire [7:0] io_out_bits_union;
	reg [31:0] data_0;
	reg [31:0] data_1;
	reg [31:0] data_2;
	reg [31:0] data_3;
	reg receiving;
	wire _T = io_in_ready & io_in_valid;
	reg [1:0] recvCount;
	wire wrap_wrap = recvCount == 2'h3;
	wire [1:0] _wrap_value_T_1 = recvCount + 2'h1;
	wire recvDone = _T & wrap_wrap;
	wire [127:0] _io_out_bits_T = {data_3, data_2, data_1, data_0};
	wire _GEN_10 = (recvDone ? 1'h0 : receiving);
	wire _T_2 = io_out_ready & io_out_valid;
	wire _GEN_11 = _T_2 | _GEN_10;
	assign io_in_ready = receiving;
	assign io_out_valid = ~receiving;
	assign io_out_bits_chanId = _io_out_bits_T[121:119];
	assign io_out_bits_opcode = _io_out_bits_T[118:116];
	assign io_out_bits_param = _io_out_bits_T[115:113];
	assign io_out_bits_size = _io_out_bits_T[112:109];
	assign io_out_bits_source = _io_out_bits_T[108:106];
	assign io_out_bits_address = _io_out_bits_T[105:74];
	assign io_out_bits_data = _io_out_bits_T[73:10];
	assign io_out_bits_corrupt = _io_out_bits_T[9];
	assign io_out_bits_union = _io_out_bits_T[8:1];
	always @(posedge clock) begin
		if (_T)
			if (2'h0 == recvCount)
				data_0 <= io_in_bits;
		if (_T)
			if (2'h1 == recvCount)
				data_1 <= io_in_bits;
		if (_T)
			if (2'h2 == recvCount)
				data_2 <= io_in_bits;
		if (_T)
			if (2'h3 == recvCount)
				data_3 <= io_in_bits;
		receiving <= reset | _GEN_11;
		if (reset)
			recvCount <= 2'h0;
		else if (_T)
			recvCount <= _wrap_value_T_1;
	end
endmodule
module TLSerdesser (
	clock,
	reset,
	auto_manager_in_a_ready,
	auto_manager_in_a_valid,
	auto_manager_in_a_bits_opcode,
	auto_manager_in_a_bits_param,
	auto_manager_in_a_bits_size,
	auto_manager_in_a_bits_source,
	auto_manager_in_a_bits_address,
	auto_manager_in_a_bits_mask,
	auto_manager_in_a_bits_data,
	auto_manager_in_a_bits_corrupt,
	auto_manager_in_d_ready,
	auto_manager_in_d_valid,
	auto_manager_in_d_bits_opcode,
	auto_manager_in_d_bits_param,
	auto_manager_in_d_bits_size,
	auto_manager_in_d_bits_source,
	auto_manager_in_d_bits_sink,
	auto_manager_in_d_bits_denied,
	auto_manager_in_d_bits_data,
	auto_manager_in_d_bits_corrupt,
	auto_client_out_a_ready,
	auto_client_out_a_valid,
	auto_client_out_a_bits_opcode,
	auto_client_out_a_bits_param,
	auto_client_out_a_bits_size,
	auto_client_out_a_bits_source,
	auto_client_out_a_bits_address,
	auto_client_out_a_bits_mask,
	auto_client_out_a_bits_data,
	auto_client_out_a_bits_corrupt,
	auto_client_out_d_ready,
	auto_client_out_d_valid,
	auto_client_out_d_bits_opcode,
	auto_client_out_d_bits_param,
	auto_client_out_d_bits_size,
	auto_client_out_d_bits_source,
	auto_client_out_d_bits_sink,
	auto_client_out_d_bits_denied,
	auto_client_out_d_bits_data,
	auto_client_out_d_bits_corrupt,
	io_ser_in_ready,
	io_ser_in_valid,
	io_ser_in_bits,
	io_ser_out_ready,
	io_ser_out_valid,
	io_ser_out_bits
);
	input clock;
	input reset;
	output wire auto_manager_in_a_ready;
	input auto_manager_in_a_valid;
	input [2:0] auto_manager_in_a_bits_opcode;
	input [2:0] auto_manager_in_a_bits_param;
	input [2:0] auto_manager_in_a_bits_size;
	input [2:0] auto_manager_in_a_bits_source;
	input [28:0] auto_manager_in_a_bits_address;
	input [7:0] auto_manager_in_a_bits_mask;
	input [63:0] auto_manager_in_a_bits_data;
	input auto_manager_in_a_bits_corrupt;
	input auto_manager_in_d_ready;
	output wire auto_manager_in_d_valid;
	output wire [2:0] auto_manager_in_d_bits_opcode;
	output wire [1:0] auto_manager_in_d_bits_param;
	output wire [2:0] auto_manager_in_d_bits_size;
	output wire [2:0] auto_manager_in_d_bits_source;
	output wire auto_manager_in_d_bits_sink;
	output wire auto_manager_in_d_bits_denied;
	output wire [63:0] auto_manager_in_d_bits_data;
	output wire auto_manager_in_d_bits_corrupt;
	input auto_client_out_a_ready;
	output wire auto_client_out_a_valid;
	output wire [2:0] auto_client_out_a_bits_opcode;
	output wire [2:0] auto_client_out_a_bits_param;
	output wire [3:0] auto_client_out_a_bits_size;
	output wire auto_client_out_a_bits_source;
	output wire [31:0] auto_client_out_a_bits_address;
	output wire [3:0] auto_client_out_a_bits_mask;
	output wire [31:0] auto_client_out_a_bits_data;
	output wire auto_client_out_a_bits_corrupt;
	output wire auto_client_out_d_ready;
	input auto_client_out_d_valid;
	input [2:0] auto_client_out_d_bits_opcode;
	input [1:0] auto_client_out_d_bits_param;
	input [3:0] auto_client_out_d_bits_size;
	input auto_client_out_d_bits_source;
	input auto_client_out_d_bits_sink;
	input auto_client_out_d_bits_denied;
	input [31:0] auto_client_out_d_bits_data;
	input auto_client_out_d_bits_corrupt;
	output wire io_ser_in_ready;
	input io_ser_in_valid;
	input [31:0] io_ser_in_bits;
	input io_ser_out_ready;
	output wire io_ser_out_valid;
	output wire [31:0] io_ser_out_bits;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [28:0] monitor_io_in_a_bits_address;
	wire [7:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire outArb_clock;
	wire outArb_reset;
	wire outArb_io_in_1_ready;
	wire outArb_io_in_1_valid;
	wire [2:0] outArb_io_in_1_bits_opcode;
	wire [2:0] outArb_io_in_1_bits_param;
	wire [3:0] outArb_io_in_1_bits_size;
	wire [2:0] outArb_io_in_1_bits_source;
	wire [63:0] outArb_io_in_1_bits_data;
	wire outArb_io_in_1_bits_corrupt;
	wire [7:0] outArb_io_in_1_bits_union;
	wire outArb_io_in_1_bits_last;
	wire outArb_io_in_4_ready;
	wire outArb_io_in_4_valid;
	wire [2:0] outArb_io_in_4_bits_opcode;
	wire [2:0] outArb_io_in_4_bits_param;
	wire [3:0] outArb_io_in_4_bits_size;
	wire [2:0] outArb_io_in_4_bits_source;
	wire [31:0] outArb_io_in_4_bits_address;
	wire [63:0] outArb_io_in_4_bits_data;
	wire outArb_io_in_4_bits_corrupt;
	wire [7:0] outArb_io_in_4_bits_union;
	wire outArb_io_in_4_bits_last;
	wire outArb_io_out_ready;
	wire outArb_io_out_valid;
	wire [2:0] outArb_io_out_bits_chanId;
	wire [2:0] outArb_io_out_bits_opcode;
	wire [2:0] outArb_io_out_bits_param;
	wire [3:0] outArb_io_out_bits_size;
	wire [2:0] outArb_io_out_bits_source;
	wire [31:0] outArb_io_out_bits_address;
	wire [63:0] outArb_io_out_bits_data;
	wire outArb_io_out_bits_corrupt;
	wire [7:0] outArb_io_out_bits_union;
	wire outArb_io_out_bits_last;
	wire outSer_clock;
	wire outSer_reset;
	wire outSer_io_in_ready;
	wire outSer_io_in_valid;
	wire [2:0] outSer_io_in_bits_chanId;
	wire [2:0] outSer_io_in_bits_opcode;
	wire [2:0] outSer_io_in_bits_param;
	wire [3:0] outSer_io_in_bits_size;
	wire [2:0] outSer_io_in_bits_source;
	wire [31:0] outSer_io_in_bits_address;
	wire [63:0] outSer_io_in_bits_data;
	wire outSer_io_in_bits_corrupt;
	wire [7:0] outSer_io_in_bits_union;
	wire outSer_io_in_bits_last;
	wire outSer_io_out_ready;
	wire outSer_io_out_valid;
	wire [31:0] outSer_io_out_bits;
	wire inDes_clock;
	wire inDes_reset;
	wire inDes_io_in_ready;
	wire inDes_io_in_valid;
	wire [31:0] inDes_io_in_bits;
	wire inDes_io_out_ready;
	wire inDes_io_out_valid;
	wire [2:0] inDes_io_out_bits_chanId;
	wire [2:0] inDes_io_out_bits_opcode;
	wire [2:0] inDes_io_out_bits_param;
	wire [3:0] inDes_io_out_bits_size;
	wire [2:0] inDes_io_out_bits_source;
	wire [31:0] inDes_io_out_bits_address;
	wire [63:0] inDes_io_out_bits_data;
	wire inDes_io_out_bits_corrupt;
	wire [7:0] inDes_io_out_bits_union;
	wire [1:0] _merged_bits_merged_union_T_1 = {auto_client_out_d_bits_sink, auto_client_out_d_bits_denied};
	wire merged_1_ready = outArb_io_in_1_ready;
	wire _merged_bits_last_T_1 = merged_1_ready & auto_client_out_d_valid;
	wire [26:0] _merged_bits_last_beats1_decode_T_1 = 27'h0000fff << auto_client_out_d_bits_size;
	wire [11:0] _merged_bits_last_beats1_decode_T_3 = ~_merged_bits_last_beats1_decode_T_1[11:0];
	wire [9:0] merged_bits_last_beats1_decode = _merged_bits_last_beats1_decode_T_3[11:2];
	wire merged_bits_last_beats1_opdata = auto_client_out_d_bits_opcode[0];
	wire [9:0] merged_bits_last_beats1 = (merged_bits_last_beats1_opdata ? merged_bits_last_beats1_decode : 10'h000);
	reg [9:0] merged_bits_last_counter_1;
	wire [9:0] merged_bits_last_counter1_1 = merged_bits_last_counter_1 - 10'h001;
	wire merged_bits_last_first_1 = merged_bits_last_counter_1 == 10'h000;
	wire merged_4_ready = outArb_io_in_4_ready;
	wire _merged_bits_last_T_4 = merged_4_ready & auto_manager_in_a_valid;
	wire [18:0] _merged_bits_last_beats1_decode_T_13 = 19'h00fff << auto_manager_in_a_bits_size;
	wire [11:0] _merged_bits_last_beats1_decode_T_15 = ~_merged_bits_last_beats1_decode_T_13[11:0];
	wire [9:0] merged_bits_last_beats1_decode_3 = _merged_bits_last_beats1_decode_T_15[11:2];
	wire merged_bits_last_beats1_opdata_3 = ~auto_manager_in_a_bits_opcode[2];
	wire [9:0] merged_bits_last_beats1_3 = (merged_bits_last_beats1_opdata_3 ? merged_bits_last_beats1_decode_3 : 10'h000);
	reg [9:0] merged_bits_last_counter_4;
	wire [9:0] merged_bits_last_counter1_4 = merged_bits_last_counter_4 - 10'h001;
	wire merged_bits_last_first_4 = merged_bits_last_counter_4 == 10'h000;
	wire _bundleOut_0_a_valid_T = inDes_io_out_bits_chanId == 3'h0;
	wire _bundleIn_0_d_valid_T = inDes_io_out_bits_chanId == 3'h3;
	wire [7:0] _bundleIn_0_d_bits_d_sink_T = {1'd0, inDes_io_out_bits_union[7:1]};
	wire _inDes_io_out_ready_T_3 = (3'h1 == inDes_io_out_bits_chanId ? 1'h0 : (3'h0 == inDes_io_out_bits_chanId) & auto_client_out_a_ready);
	wire _inDes_io_out_ready_T_5 = (3'h2 == inDes_io_out_bits_chanId ? 1'h0 : _inDes_io_out_ready_T_3);
	wire _inDes_io_out_ready_T_7 = (3'h3 == inDes_io_out_bits_chanId ? auto_manager_in_d_ready : _inDes_io_out_ready_T_5);
	TLMonitor_44 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	HellaPeekingArbiter outArb(
		.clock(outArb_clock),
		.reset(outArb_reset),
		.io_in_1_ready(outArb_io_in_1_ready),
		.io_in_1_valid(outArb_io_in_1_valid),
		.io_in_1_bits_opcode(outArb_io_in_1_bits_opcode),
		.io_in_1_bits_param(outArb_io_in_1_bits_param),
		.io_in_1_bits_size(outArb_io_in_1_bits_size),
		.io_in_1_bits_source(outArb_io_in_1_bits_source),
		.io_in_1_bits_data(outArb_io_in_1_bits_data),
		.io_in_1_bits_corrupt(outArb_io_in_1_bits_corrupt),
		.io_in_1_bits_union(outArb_io_in_1_bits_union),
		.io_in_1_bits_last(outArb_io_in_1_bits_last),
		.io_in_4_ready(outArb_io_in_4_ready),
		.io_in_4_valid(outArb_io_in_4_valid),
		.io_in_4_bits_opcode(outArb_io_in_4_bits_opcode),
		.io_in_4_bits_param(outArb_io_in_4_bits_param),
		.io_in_4_bits_size(outArb_io_in_4_bits_size),
		.io_in_4_bits_source(outArb_io_in_4_bits_source),
		.io_in_4_bits_address(outArb_io_in_4_bits_address),
		.io_in_4_bits_data(outArb_io_in_4_bits_data),
		.io_in_4_bits_corrupt(outArb_io_in_4_bits_corrupt),
		.io_in_4_bits_union(outArb_io_in_4_bits_union),
		.io_in_4_bits_last(outArb_io_in_4_bits_last),
		.io_out_ready(outArb_io_out_ready),
		.io_out_valid(outArb_io_out_valid),
		.io_out_bits_chanId(outArb_io_out_bits_chanId),
		.io_out_bits_opcode(outArb_io_out_bits_opcode),
		.io_out_bits_param(outArb_io_out_bits_param),
		.io_out_bits_size(outArb_io_out_bits_size),
		.io_out_bits_source(outArb_io_out_bits_source),
		.io_out_bits_address(outArb_io_out_bits_address),
		.io_out_bits_data(outArb_io_out_bits_data),
		.io_out_bits_corrupt(outArb_io_out_bits_corrupt),
		.io_out_bits_union(outArb_io_out_bits_union),
		.io_out_bits_last(outArb_io_out_bits_last)
	);
	GenericSerializer outSer(
		.clock(outSer_clock),
		.reset(outSer_reset),
		.io_in_ready(outSer_io_in_ready),
		.io_in_valid(outSer_io_in_valid),
		.io_in_bits_chanId(outSer_io_in_bits_chanId),
		.io_in_bits_opcode(outSer_io_in_bits_opcode),
		.io_in_bits_param(outSer_io_in_bits_param),
		.io_in_bits_size(outSer_io_in_bits_size),
		.io_in_bits_source(outSer_io_in_bits_source),
		.io_in_bits_address(outSer_io_in_bits_address),
		.io_in_bits_data(outSer_io_in_bits_data),
		.io_in_bits_corrupt(outSer_io_in_bits_corrupt),
		.io_in_bits_union(outSer_io_in_bits_union),
		.io_in_bits_last(outSer_io_in_bits_last),
		.io_out_ready(outSer_io_out_ready),
		.io_out_valid(outSer_io_out_valid),
		.io_out_bits(outSer_io_out_bits)
	);
	GenericDeserializer inDes(
		.clock(inDes_clock),
		.reset(inDes_reset),
		.io_in_ready(inDes_io_in_ready),
		.io_in_valid(inDes_io_in_valid),
		.io_in_bits(inDes_io_in_bits),
		.io_out_ready(inDes_io_out_ready),
		.io_out_valid(inDes_io_out_valid),
		.io_out_bits_chanId(inDes_io_out_bits_chanId),
		.io_out_bits_opcode(inDes_io_out_bits_opcode),
		.io_out_bits_param(inDes_io_out_bits_param),
		.io_out_bits_size(inDes_io_out_bits_size),
		.io_out_bits_source(inDes_io_out_bits_source),
		.io_out_bits_address(inDes_io_out_bits_address),
		.io_out_bits_data(inDes_io_out_bits_data),
		.io_out_bits_corrupt(inDes_io_out_bits_corrupt),
		.io_out_bits_union(inDes_io_out_bits_union)
	);
	assign auto_manager_in_a_ready = outArb_io_in_4_ready;
	assign auto_manager_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T;
	assign auto_manager_in_d_bits_opcode = inDes_io_out_bits_opcode;
	assign auto_manager_in_d_bits_param = inDes_io_out_bits_param[1:0];
	assign auto_manager_in_d_bits_size = inDes_io_out_bits_size[2:0];
	assign auto_manager_in_d_bits_source = inDes_io_out_bits_source;
	assign auto_manager_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[0];
	assign auto_manager_in_d_bits_denied = inDes_io_out_bits_union[0];
	assign auto_manager_in_d_bits_data = inDes_io_out_bits_data;
	assign auto_manager_in_d_bits_corrupt = inDes_io_out_bits_corrupt;
	assign auto_client_out_a_valid = inDes_io_out_valid & _bundleOut_0_a_valid_T;
	assign auto_client_out_a_bits_opcode = inDes_io_out_bits_opcode;
	assign auto_client_out_a_bits_param = inDes_io_out_bits_param;
	assign auto_client_out_a_bits_size = inDes_io_out_bits_size;
	assign auto_client_out_a_bits_source = inDes_io_out_bits_source[0];
	assign auto_client_out_a_bits_address = inDes_io_out_bits_address;
	assign auto_client_out_a_bits_mask = inDes_io_out_bits_union[3:0];
	assign auto_client_out_a_bits_data = inDes_io_out_bits_data[31:0];
	assign auto_client_out_a_bits_corrupt = inDes_io_out_bits_corrupt;
	assign auto_client_out_d_ready = outArb_io_in_1_ready;
	assign io_ser_in_ready = inDes_io_in_ready;
	assign io_ser_out_valid = outSer_io_out_valid;
	assign io_ser_out_bits = outSer_io_out_bits;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = outArb_io_in_4_ready;
	assign monitor_io_in_a_valid = auto_manager_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_manager_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_manager_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_manager_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_manager_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_manager_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_manager_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_manager_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_manager_in_d_ready;
	assign monitor_io_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T;
	assign monitor_io_in_d_bits_opcode = inDes_io_out_bits_opcode;
	assign monitor_io_in_d_bits_param = inDes_io_out_bits_param[1:0];
	assign monitor_io_in_d_bits_size = inDes_io_out_bits_size[2:0];
	assign monitor_io_in_d_bits_source = inDes_io_out_bits_source;
	assign monitor_io_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[0];
	assign monitor_io_in_d_bits_denied = inDes_io_out_bits_union[0];
	assign monitor_io_in_d_bits_corrupt = inDes_io_out_bits_corrupt;
	assign outArb_clock = clock;
	assign outArb_reset = reset;
	assign outArb_io_in_1_valid = auto_client_out_d_valid;
	assign outArb_io_in_1_bits_opcode = auto_client_out_d_bits_opcode;
	assign outArb_io_in_1_bits_param = {1'd0, auto_client_out_d_bits_param};
	assign outArb_io_in_1_bits_size = auto_client_out_d_bits_size;
	assign outArb_io_in_1_bits_source = {2'd0, auto_client_out_d_bits_source};
	assign outArb_io_in_1_bits_data = {32'd0, auto_client_out_d_bits_data};
	assign outArb_io_in_1_bits_corrupt = auto_client_out_d_bits_corrupt;
	assign outArb_io_in_1_bits_union = {6'd0, _merged_bits_merged_union_T_1};
	assign outArb_io_in_1_bits_last = (merged_bits_last_counter_1 == 10'h001) | (merged_bits_last_beats1 == 10'h000);
	assign outArb_io_in_4_valid = auto_manager_in_a_valid;
	assign outArb_io_in_4_bits_opcode = auto_manager_in_a_bits_opcode;
	assign outArb_io_in_4_bits_param = auto_manager_in_a_bits_param;
	assign outArb_io_in_4_bits_size = {1'd0, auto_manager_in_a_bits_size};
	assign outArb_io_in_4_bits_source = auto_manager_in_a_bits_source;
	assign outArb_io_in_4_bits_address = {3'd0, auto_manager_in_a_bits_address};
	assign outArb_io_in_4_bits_data = auto_manager_in_a_bits_data;
	assign outArb_io_in_4_bits_corrupt = auto_manager_in_a_bits_corrupt;
	assign outArb_io_in_4_bits_union = auto_manager_in_a_bits_mask;
	assign outArb_io_in_4_bits_last = (merged_bits_last_counter_4 == 10'h001) | (merged_bits_last_beats1_3 == 10'h000);
	assign outArb_io_out_ready = outSer_io_in_ready;
	assign outSer_clock = clock;
	assign outSer_reset = reset;
	assign outSer_io_in_valid = outArb_io_out_valid;
	assign outSer_io_in_bits_chanId = outArb_io_out_bits_chanId;
	assign outSer_io_in_bits_opcode = outArb_io_out_bits_opcode;
	assign outSer_io_in_bits_param = outArb_io_out_bits_param;
	assign outSer_io_in_bits_size = outArb_io_out_bits_size;
	assign outSer_io_in_bits_source = outArb_io_out_bits_source;
	assign outSer_io_in_bits_address = outArb_io_out_bits_address;
	assign outSer_io_in_bits_data = outArb_io_out_bits_data;
	assign outSer_io_in_bits_corrupt = outArb_io_out_bits_corrupt;
	assign outSer_io_in_bits_union = outArb_io_out_bits_union;
	assign outSer_io_in_bits_last = outArb_io_out_bits_last;
	assign outSer_io_out_ready = io_ser_out_ready;
	assign inDes_clock = clock;
	assign inDes_reset = reset;
	assign inDes_io_in_valid = io_ser_in_valid;
	assign inDes_io_in_bits = io_ser_in_bits;
	assign inDes_io_out_ready = (3'h4 == inDes_io_out_bits_chanId ? 1'h0 : _inDes_io_out_ready_T_7);
	always @(posedge clock) begin
		if (reset)
			merged_bits_last_counter_1 <= 10'h000;
		else if (_merged_bits_last_T_1)
			if (merged_bits_last_first_1) begin
				if (merged_bits_last_beats1_opdata)
					merged_bits_last_counter_1 <= merged_bits_last_beats1_decode;
				else
					merged_bits_last_counter_1 <= 10'h000;
			end
			else
				merged_bits_last_counter_1 <= merged_bits_last_counter1_1;
		if (reset)
			merged_bits_last_counter_4 <= 10'h000;
		else if (_merged_bits_last_T_4)
			if (merged_bits_last_first_4) begin
				if (merged_bits_last_beats1_opdata_3)
					merged_bits_last_counter_4 <= merged_bits_last_beats1_decode_3;
				else
					merged_bits_last_counter_4 <= 10'h000;
			end
			else
				merged_bits_last_counter_4 <= merged_bits_last_counter1_4;
	end
endmodule
module TLMonitor_45 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [2:0] io_in_a_bits_size;
	input [2:0] io_in_a_bits_source;
	input [28:0] io_in_a_bits_address;
	input [7:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [2:0] io_in_d_bits_size;
	input [2:0] io_in_d_bits_source;
	input io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T = io_in_a_bits_source == 3'h2;
	wire _source_ok_T_1 = io_in_a_bits_source == 3'h1;
	wire _source_ok_T_2 = io_in_a_bits_source == 3'h0;
	wire _source_ok_T_3 = io_in_a_bits_source == 3'h4;
	wire source_ok = ((_source_ok_T | _source_ok_T_1) | _source_ok_T_2) | _source_ok_T_3;
	wire [12:0] _is_aligned_mask_T_1 = 13'h003f << io_in_a_bits_size;
	wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0];
	wire [28:0] _GEN_71 = {23'd0, is_aligned_mask};
	wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 29'h00000000;
	wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0];
	wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount;
	wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1;
	wire _mask_T = io_in_a_bits_size >= 3'h3;
	wire mask_size = mask_sizeOH[2];
	wire mask_bit = io_in_a_bits_address[2];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[1];
	wire mask_bit_1 = io_in_a_bits_address[1];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire mask_size_2 = mask_sizeOH[0];
	wire mask_bit_2 = io_in_a_bits_address[0];
	wire mask_nbit_2 = ~mask_bit_2;
	wire mask_eq_6 = mask_eq_2 & mask_nbit_2;
	wire mask_acc_6 = mask_acc_2 | (mask_size_2 & mask_eq_6);
	wire mask_eq_7 = mask_eq_2 & mask_bit_2;
	wire mask_acc_7 = mask_acc_2 | (mask_size_2 & mask_eq_7);
	wire mask_eq_8 = mask_eq_3 & mask_nbit_2;
	wire mask_acc_8 = mask_acc_3 | (mask_size_2 & mask_eq_8);
	wire mask_eq_9 = mask_eq_3 & mask_bit_2;
	wire mask_acc_9 = mask_acc_3 | (mask_size_2 & mask_eq_9);
	wire mask_eq_10 = mask_eq_4 & mask_nbit_2;
	wire mask_acc_10 = mask_acc_4 | (mask_size_2 & mask_eq_10);
	wire mask_eq_11 = mask_eq_4 & mask_bit_2;
	wire mask_acc_11 = mask_acc_4 | (mask_size_2 & mask_eq_11);
	wire mask_eq_12 = mask_eq_5 & mask_nbit_2;
	wire mask_acc_12 = mask_acc_5 | (mask_size_2 & mask_eq_12);
	wire mask_eq_13 = mask_eq_5 & mask_bit_2;
	wire mask_acc_13 = mask_acc_5 | (mask_size_2 & mask_eq_13);
	wire [7:0] mask = {mask_acc_13, mask_acc_12, mask_acc_11, mask_acc_10, mask_acc_9, mask_acc_8, mask_acc_7, mask_acc_6};
	wire _T_42 = io_in_a_bits_opcode == 3'h6;
	wire [28:0] _T_56 = io_in_a_bits_address ^ 29'h00020000;
	wire [29:0] _T_57 = {1'b0, $signed(_T_56)};
	wire [29:0] _T_59 = $signed(_T_57) & -30'sh00010000;
	wire _T_60 = $signed(_T_59) == 30'sh00000000;
	wire [28:0] _T_61 = io_in_a_bits_address ^ 29'h10000000;
	wire [29:0] _T_62 = {1'b0, $signed(_T_61)};
	wire [29:0] _T_64 = $signed(_T_62) & -30'sh00001000;
	wire _T_65 = $signed(_T_64) == 30'sh00000000;
	wire _T_66 = _T_60 | _T_65;
	wire _T_104 = io_in_a_bits_param <= 3'h2;
	wire [7:0] _T_108 = ~io_in_a_bits_mask;
	wire _T_109 = _T_108 == 8'h00;
	wire _T_113 = ~io_in_a_bits_corrupt;
	wire _T_117 = io_in_a_bits_opcode == 3'h7;
	wire _T_183 = io_in_a_bits_param != 3'h0;
	wire _T_196 = io_in_a_bits_opcode == 3'h4;
	wire _T_213 = io_in_a_bits_size <= 3'h6;
	wire _T_227 = _T_213 & _T_66;
	wire _T_238 = io_in_a_bits_param == 3'h0;
	wire _T_242 = io_in_a_bits_mask == mask;
	wire _T_250 = io_in_a_bits_opcode == 3'h0;
	wire _T_272 = _T_213 & _T_65;
	wire _T_282 = source_ok & _T_272;
	wire _T_300 = io_in_a_bits_opcode == 3'h1;
	wire [7:0] _T_346 = ~mask;
	wire [7:0] _T_347 = io_in_a_bits_mask & _T_346;
	wire _T_348 = _T_347 == 8'h00;
	wire _T_352 = io_in_a_bits_opcode == 3'h2;
	wire _T_389 = io_in_a_bits_param <= 3'h4;
	wire _T_397 = io_in_a_bits_opcode == 3'h3;
	wire _T_434 = io_in_a_bits_param <= 3'h3;
	wire _T_442 = io_in_a_bits_opcode == 3'h5;
	wire _T_479 = io_in_a_bits_param <= 3'h1;
	wire _T_491 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_6 = io_in_d_bits_source == 3'h2;
	wire _source_ok_T_7 = io_in_d_bits_source == 3'h1;
	wire _source_ok_T_8 = io_in_d_bits_source == 3'h0;
	wire _source_ok_T_9 = io_in_d_bits_source == 3'h4;
	wire source_ok_1 = ((_source_ok_T_6 | _source_ok_T_7) | _source_ok_T_8) | _source_ok_T_9;
	wire _T_495 = io_in_d_bits_opcode == 3'h6;
	wire _T_499 = io_in_d_bits_size >= 3'h3;
	wire _T_503 = io_in_d_bits_param == 2'h0;
	wire _T_507 = ~io_in_d_bits_corrupt;
	wire _T_511 = ~io_in_d_bits_denied;
	wire _T_515 = io_in_d_bits_opcode == 3'h4;
	wire _T_526 = io_in_d_bits_param <= 2'h2;
	wire _T_530 = io_in_d_bits_param != 2'h2;
	wire _T_543 = io_in_d_bits_opcode == 3'h5;
	wire _T_563 = _T_511 | io_in_d_bits_corrupt;
	wire _T_572 = io_in_d_bits_opcode == 3'h0;
	wire _T_589 = io_in_d_bits_opcode == 3'h1;
	wire _T_607 = io_in_d_bits_opcode == 3'h2;
	wire _a_first_T = io_in_a_ready & io_in_a_valid;
	wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3];
	wire a_first_beats1_opdata = ~io_in_a_bits_opcode[2];
	reg [2:0] a_first_counter;
	wire [2:0] a_first_counter1 = a_first_counter - 3'h1;
	wire a_first = a_first_counter == 3'h0;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [2:0] size;
	reg [2:0] source;
	reg [28:0] address;
	wire _T_637 = io_in_a_valid & ~a_first;
	wire _T_638 = io_in_a_bits_opcode == opcode;
	wire _T_642 = io_in_a_bits_param == param;
	wire _T_646 = io_in_a_bits_size == size;
	wire _T_650 = io_in_a_bits_source == source;
	wire _T_654 = io_in_a_bits_address == address;
	wire _d_first_T = io_in_d_ready & io_in_d_valid;
	wire [12:0] _d_first_beats1_decode_T_1 = 13'h003f << io_in_d_bits_size;
	wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0];
	wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3];
	wire d_first_beats1_opdata = io_in_d_bits_opcode[0];
	reg [2:0] d_first_counter;
	wire [2:0] d_first_counter1 = d_first_counter - 3'h1;
	wire d_first = d_first_counter == 3'h0;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [2:0] size_1;
	reg [2:0] source_1;
	reg sink;
	reg denied;
	wire _T_661 = io_in_d_valid & ~d_first;
	wire _T_662 = io_in_d_bits_opcode == opcode_1;
	wire _T_666 = io_in_d_bits_param == param_1;
	wire _T_670 = io_in_d_bits_size == size_1;
	wire _T_674 = io_in_d_bits_source == source_1;
	wire _T_678 = io_in_d_bits_sink == sink;
	wire _T_682 = io_in_d_bits_denied == denied;
	reg [4:0] inflight;
	reg [19:0] inflight_opcodes;
	reg [19:0] inflight_sizes;
	reg [2:0] a_first_counter_1;
	wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1;
	wire a_first_1 = a_first_counter_1 == 3'h0;
	reg [2:0] d_first_counter_1;
	wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1;
	wire d_first_1 = d_first_counter_1 == 3'h0;
	wire [4:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [5:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [19:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [19:0] _GEN_73 = {4'd0, _a_opcode_lookup_T_5};
	wire [19:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [19:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[19:1]};
	wire [19:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [19:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [19:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[19:1]};
	wire _T_688 = io_in_a_valid & a_first_1;
	wire [7:0] _a_set_wo_ready_T = 8'h01 << io_in_a_bits_source;
	wire [7:0] _GEN_15 = (io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire _T_691 = _a_first_T & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1;
	wire [4:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [5:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (_a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_1 = {63'd0, a_opcodes_set_interm};
	wire [66:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [3:0] a_sizes_set_interm = (_a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0);
	wire [66:0] _GEN_2 = {63'd0, a_sizes_set_interm};
	wire [66:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [4:0] _T_693 = inflight >> io_in_a_bits_source;
	wire _T_695 = ~_T_693[0];
	wire [7:0] _GEN_16 = (_a_first_T & a_first_1 ? _a_set_wo_ready_T : 8'h00);
	wire [66:0] _GEN_19 = (_a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 67'h00000000000000000);
	wire [66:0] _GEN_20 = (_a_first_T & a_first_1 ? _a_sizes_set_T_1 : 67'h00000000000000000);
	wire _T_699 = io_in_d_valid & d_first_1;
	wire _T_701 = ~_T_495;
	wire _T_702 = (io_in_d_valid & d_first_1) & ~_T_495;
	wire [7:0] _d_clr_wo_ready_T = 8'h01 << io_in_d_bits_source;
	wire [7:0] _GEN_21 = ((io_in_d_valid & d_first_1) & ~_T_495 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_3 = {63'd0, _a_opcode_lookup_T_5};
	wire [78:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [7:0] _GEN_22 = ((_d_first_T & d_first_1) & _T_701 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_23 = ((_d_first_T & d_first_1) & _T_701 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_688 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [4:0] _T_712 = inflight >> io_in_d_bits_source;
	wire _T_714 = _T_712[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_719 = io_in_d_bits_opcode == _GEN_40;
	wire _T_720 = (io_in_d_bits_opcode == _GEN_32) | _T_719;
	wire _T_724 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_731 = io_in_d_bits_opcode == _GEN_56;
	wire _T_732 = (io_in_d_bits_opcode == _GEN_48) | _T_731;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {1'd0, io_in_d_bits_size};
	wire _T_736 = _GEN_82 == a_size_lookup;
	wire _T_746 = (((_T_699 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_701;
	wire _T_748 = ~io_in_d_ready | io_in_a_ready;
	wire [4:0] a_set_wo_ready = _GEN_15[4:0];
	wire [4:0] d_clr_wo_ready = _GEN_21[4:0];
	wire _T_755 = (a_set_wo_ready != d_clr_wo_ready) | ~(|a_set_wo_ready);
	wire [4:0] a_set = _GEN_16[4:0];
	wire [4:0] _inflight_T = inflight | a_set;
	wire [4:0] d_clr = _GEN_22[4:0];
	wire [4:0] _inflight_T_1 = ~d_clr;
	wire [4:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [19:0] a_opcodes_set = _GEN_19[19:0];
	wire [19:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [19:0] d_opcodes_clr = _GEN_23[19:0];
	wire [19:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [19:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [19:0] a_sizes_set = _GEN_20[19:0];
	wire [19:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [19:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_764 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [4:0] inflight_1;
	reg [19:0] inflight_sizes_1;
	reg [2:0] d_first_counter_2;
	wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1;
	wire d_first_2 = d_first_counter_2 == 3'h0;
	wire [19:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [19:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [19:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[19:1]};
	wire _T_790 = (io_in_d_valid & d_first_2) & _T_495;
	wire [7:0] _GEN_67 = ((_d_first_T & d_first_2) & _T_495 ? _d_clr_wo_ready_T : 8'h00);
	wire [78:0] _GEN_68 = ((_d_first_T & d_first_2) & _T_495 ? _d_opcodes_clr_T_5 : 79'h00000000000000000000);
	wire [4:0] _T_798 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_808 = _GEN_82 == c_size_lookup;
	wire [4:0] d_clr_1 = _GEN_67[4:0];
	wire [4:0] _inflight_T_4 = ~d_clr_1;
	wire [4:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [19:0] d_opcodes_clr_1 = _GEN_68[19:0];
	wire [19:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [19:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_833 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 3'h0;
		else if (_a_first_T)
			if (a_first) begin
				if (a_first_beats1_opdata)
					a_first_counter <= a_first_beats1_decode;
				else
					a_first_counter <= 3'h0;
			end
			else
				a_first_counter <= a_first_counter1;
		if (_a_first_T & a_first)
			opcode <= io_in_a_bits_opcode;
		if (_a_first_T & a_first)
			param <= io_in_a_bits_param;
		if (_a_first_T & a_first)
			size <= io_in_a_bits_size;
		if (_a_first_T & a_first)
			source <= io_in_a_bits_source;
		if (_a_first_T & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 3'h0;
		else if (_d_first_T)
			if (d_first) begin
				if (d_first_beats1_opdata)
					d_first_counter <= d_first_beats1_decode;
				else
					d_first_counter <= 3'h0;
			end
			else
				d_first_counter <= d_first_counter1;
		if (_d_first_T & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (_d_first_T & d_first)
			param_1 <= io_in_d_bits_param;
		if (_d_first_T & d_first)
			size_1 <= io_in_d_bits_size;
		if (_d_first_T & d_first)
			source_1 <= io_in_d_bits_source;
		if (_d_first_T & d_first)
			sink <= io_in_d_bits_sink;
		if (_d_first_T & d_first)
			denied <= io_in_d_bits_denied;
		if (reset)
			inflight <= 5'h00;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 20'h00000;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 20'h00000;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 3'h0;
		else if (_a_first_T)
			if (a_first_1) begin
				if (a_first_beats1_opdata)
					a_first_counter_1 <= a_first_beats1_decode;
				else
					a_first_counter_1 <= 3'h0;
			end
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 3'h0;
		else if (_d_first_T)
			if (d_first_1) begin
				if (d_first_beats1_opdata)
					d_first_counter_1 <= d_first_beats1_decode;
				else
					d_first_counter_1 <= 3'h0;
			end
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (_a_first_T | _d_first_T)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 5'h00;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 20'h00000;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 3'h0;
		else if (_d_first_T)
			if (d_first_2) begin
				if (d_first_beats1_opdata)
					d_first_counter_2 <= d_first_beats1_decode;
				else
					d_first_counter_2 <= 3'h0;
			end
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (_d_first_T)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module Queue_22 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_data,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input [28:0] io_enq_bits_address;
	input [7:0] io_enq_bits_mask;
	input [63:0] io_enq_bits_data;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire [28:0] io_deq_bits_address;
	output wire [7:0] io_deq_bits_mask;
	output wire [63:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg [2:0] ram_opcode [0:1];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [2:0] ram_param [0:1];
	wire ram_param_io_deq_bits_MPORT_en;
	wire ram_param_io_deq_bits_MPORT_addr;
	wire [2:0] ram_param_io_deq_bits_MPORT_data;
	wire [2:0] ram_param_MPORT_data;
	wire ram_param_MPORT_addr;
	wire ram_param_MPORT_mask;
	wire ram_param_MPORT_en;
	reg [2:0] ram_size [0:1];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [2:0] ram_size_io_deq_bits_MPORT_data;
	wire [2:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg [2:0] ram_source [0:1];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire [2:0] ram_source_io_deq_bits_MPORT_data;
	wire [2:0] ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg [28:0] ram_address [0:1];
	wire ram_address_io_deq_bits_MPORT_en;
	wire ram_address_io_deq_bits_MPORT_addr;
	wire [28:0] ram_address_io_deq_bits_MPORT_data;
	wire [28:0] ram_address_MPORT_data;
	wire ram_address_MPORT_addr;
	wire ram_address_MPORT_mask;
	wire ram_address_MPORT_en;
	reg [7:0] ram_mask [0:1];
	wire ram_mask_io_deq_bits_MPORT_en;
	wire ram_mask_io_deq_bits_MPORT_addr;
	wire [7:0] ram_mask_io_deq_bits_MPORT_data;
	wire [7:0] ram_mask_MPORT_data;
	wire ram_mask_MPORT_addr;
	wire ram_mask_MPORT_mask;
	wire ram_mask_MPORT_en;
	reg [63:0] ram_data [0:1];
	wire ram_data_io_deq_bits_MPORT_en;
	wire ram_data_io_deq_bits_MPORT_addr;
	wire [63:0] ram_data_io_deq_bits_MPORT_data;
	wire [63:0] ram_data_MPORT_data;
	wire ram_data_MPORT_addr;
	wire ram_data_MPORT_mask;
	wire ram_data_MPORT_en;
	reg ram_corrupt [0:1];
	wire ram_corrupt_io_deq_bits_MPORT_en;
	wire ram_corrupt_io_deq_bits_MPORT_addr;
	wire ram_corrupt_io_deq_bits_MPORT_data;
	wire ram_corrupt_MPORT_data;
	wire ram_corrupt_MPORT_addr;
	wire ram_corrupt_MPORT_mask;
	wire ram_corrupt_MPORT_en;
	reg value;
	reg value_1;
	reg maybe_full;
	wire ptr_match = value == value_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = value;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_param_io_deq_bits_MPORT_en = 1'h1;
	assign ram_param_io_deq_bits_MPORT_addr = value_1;
	assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr];
	assign ram_param_MPORT_data = io_enq_bits_param;
	assign ram_param_MPORT_addr = value;
	assign ram_param_MPORT_mask = 1'h1;
	assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = value_1;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = value;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = value_1;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = value;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_address_io_deq_bits_MPORT_en = 1'h1;
	assign ram_address_io_deq_bits_MPORT_addr = value_1;
	assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr];
	assign ram_address_MPORT_data = io_enq_bits_address;
	assign ram_address_MPORT_addr = value;
	assign ram_address_MPORT_mask = 1'h1;
	assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
	assign ram_mask_io_deq_bits_MPORT_addr = value_1;
	assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr];
	assign ram_mask_MPORT_data = io_enq_bits_mask;
	assign ram_mask_MPORT_addr = value;
	assign ram_mask_MPORT_mask = 1'h1;
	assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_data_io_deq_bits_MPORT_en = 1'h1;
	assign ram_data_io_deq_bits_MPORT_addr = value_1;
	assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr];
	assign ram_data_MPORT_data = io_enq_bits_data;
	assign ram_data_MPORT_addr = value;
	assign ram_data_MPORT_mask = 1'h1;
	assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
	assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
	assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr];
	assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
	assign ram_corrupt_MPORT_addr = value;
	assign ram_corrupt_MPORT_mask = 1'h1;
	assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data;
	assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data;
	assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data;
	assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_param_MPORT_en & ram_param_MPORT_mask)
			ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (ram_address_MPORT_en & ram_address_MPORT_mask)
			ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data;
		if (ram_mask_MPORT_en & ram_mask_MPORT_mask)
			ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data;
		if (ram_data_MPORT_en & ram_data_MPORT_mask)
			ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data;
		if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask)
			ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data;
		if (reset)
			value <= 1'h0;
		else if (do_enq)
			value <= value + 1'h1;
		if (reset)
			value_1 <= 1'h0;
		else if (do_deq)
			value_1 <= value_1 + 1'h1;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module Queue_23 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_sink,
	io_enq_bits_denied,
	io_enq_bits_data,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_sink,
	io_deq_bits_denied,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [1:0] io_enq_bits_param;
	input [2:0] io_enq_bits_size;
	input [2:0] io_enq_bits_source;
	input io_enq_bits_sink;
	input io_enq_bits_denied;
	input [63:0] io_enq_bits_data;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [1:0] io_deq_bits_param;
	output wire [2:0] io_deq_bits_size;
	output wire [2:0] io_deq_bits_source;
	output wire io_deq_bits_sink;
	output wire io_deq_bits_denied;
	output wire [63:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg [2:0] ram_opcode [0:1];
	wire ram_opcode_io_deq_bits_MPORT_en;
	wire ram_opcode_io_deq_bits_MPORT_addr;
	wire [2:0] ram_opcode_io_deq_bits_MPORT_data;
	wire [2:0] ram_opcode_MPORT_data;
	wire ram_opcode_MPORT_addr;
	wire ram_opcode_MPORT_mask;
	wire ram_opcode_MPORT_en;
	reg [1:0] ram_param [0:1];
	wire ram_param_io_deq_bits_MPORT_en;
	wire ram_param_io_deq_bits_MPORT_addr;
	wire [1:0] ram_param_io_deq_bits_MPORT_data;
	wire [1:0] ram_param_MPORT_data;
	wire ram_param_MPORT_addr;
	wire ram_param_MPORT_mask;
	wire ram_param_MPORT_en;
	reg [2:0] ram_size [0:1];
	wire ram_size_io_deq_bits_MPORT_en;
	wire ram_size_io_deq_bits_MPORT_addr;
	wire [2:0] ram_size_io_deq_bits_MPORT_data;
	wire [2:0] ram_size_MPORT_data;
	wire ram_size_MPORT_addr;
	wire ram_size_MPORT_mask;
	wire ram_size_MPORT_en;
	reg [2:0] ram_source [0:1];
	wire ram_source_io_deq_bits_MPORT_en;
	wire ram_source_io_deq_bits_MPORT_addr;
	wire [2:0] ram_source_io_deq_bits_MPORT_data;
	wire [2:0] ram_source_MPORT_data;
	wire ram_source_MPORT_addr;
	wire ram_source_MPORT_mask;
	wire ram_source_MPORT_en;
	reg ram_sink [0:1];
	wire ram_sink_io_deq_bits_MPORT_en;
	wire ram_sink_io_deq_bits_MPORT_addr;
	wire ram_sink_io_deq_bits_MPORT_data;
	wire ram_sink_MPORT_data;
	wire ram_sink_MPORT_addr;
	wire ram_sink_MPORT_mask;
	wire ram_sink_MPORT_en;
	reg ram_denied [0:1];
	wire ram_denied_io_deq_bits_MPORT_en;
	wire ram_denied_io_deq_bits_MPORT_addr;
	wire ram_denied_io_deq_bits_MPORT_data;
	wire ram_denied_MPORT_data;
	wire ram_denied_MPORT_addr;
	wire ram_denied_MPORT_mask;
	wire ram_denied_MPORT_en;
	reg [63:0] ram_data [0:1];
	wire ram_data_io_deq_bits_MPORT_en;
	wire ram_data_io_deq_bits_MPORT_addr;
	wire [63:0] ram_data_io_deq_bits_MPORT_data;
	wire [63:0] ram_data_MPORT_data;
	wire ram_data_MPORT_addr;
	wire ram_data_MPORT_mask;
	wire ram_data_MPORT_en;
	reg ram_corrupt [0:1];
	wire ram_corrupt_io_deq_bits_MPORT_en;
	wire ram_corrupt_io_deq_bits_MPORT_addr;
	wire ram_corrupt_io_deq_bits_MPORT_data;
	wire ram_corrupt_MPORT_data;
	wire ram_corrupt_MPORT_addr;
	wire ram_corrupt_MPORT_mask;
	wire ram_corrupt_MPORT_en;
	reg value;
	reg value_1;
	reg maybe_full;
	wire ptr_match = value == value_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
	assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
	assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr];
	assign ram_opcode_MPORT_data = io_enq_bits_opcode;
	assign ram_opcode_MPORT_addr = value;
	assign ram_opcode_MPORT_mask = 1'h1;
	assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_param_io_deq_bits_MPORT_en = 1'h1;
	assign ram_param_io_deq_bits_MPORT_addr = value_1;
	assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr];
	assign ram_param_MPORT_data = io_enq_bits_param;
	assign ram_param_MPORT_addr = value;
	assign ram_param_MPORT_mask = 1'h1;
	assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_size_io_deq_bits_MPORT_en = 1'h1;
	assign ram_size_io_deq_bits_MPORT_addr = value_1;
	assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr];
	assign ram_size_MPORT_data = io_enq_bits_size;
	assign ram_size_MPORT_addr = value;
	assign ram_size_MPORT_mask = 1'h1;
	assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_source_io_deq_bits_MPORT_en = 1'h1;
	assign ram_source_io_deq_bits_MPORT_addr = value_1;
	assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr];
	assign ram_source_MPORT_data = io_enq_bits_source;
	assign ram_source_MPORT_addr = value;
	assign ram_source_MPORT_mask = 1'h1;
	assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_sink_io_deq_bits_MPORT_en = 1'h1;
	assign ram_sink_io_deq_bits_MPORT_addr = value_1;
	assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr];
	assign ram_sink_MPORT_data = io_enq_bits_sink;
	assign ram_sink_MPORT_addr = value;
	assign ram_sink_MPORT_mask = 1'h1;
	assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_denied_io_deq_bits_MPORT_en = 1'h1;
	assign ram_denied_io_deq_bits_MPORT_addr = value_1;
	assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr];
	assign ram_denied_MPORT_data = io_enq_bits_denied;
	assign ram_denied_MPORT_addr = value;
	assign ram_denied_MPORT_mask = 1'h1;
	assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_data_io_deq_bits_MPORT_en = 1'h1;
	assign ram_data_io_deq_bits_MPORT_addr = value_1;
	assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr];
	assign ram_data_MPORT_data = io_enq_bits_data;
	assign ram_data_MPORT_addr = value;
	assign ram_data_MPORT_mask = 1'h1;
	assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
	assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
	assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
	assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr];
	assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
	assign ram_corrupt_MPORT_addr = value;
	assign ram_corrupt_MPORT_mask = 1'h1;
	assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data;
	assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data;
	assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data;
	assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data;
	assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data;
	assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data;
	assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data;
	assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data;
	always @(posedge clock) begin
		if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask)
			ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data;
		if (ram_param_MPORT_en & ram_param_MPORT_mask)
			ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data;
		if (ram_size_MPORT_en & ram_size_MPORT_mask)
			ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data;
		if (ram_source_MPORT_en & ram_source_MPORT_mask)
			ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data;
		if (ram_sink_MPORT_en & ram_sink_MPORT_mask)
			ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data;
		if (ram_denied_MPORT_en & ram_denied_MPORT_mask)
			ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data;
		if (ram_data_MPORT_en & ram_data_MPORT_mask)
			ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data;
		if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask)
			ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data;
		if (reset)
			value <= 1'h0;
		else if (do_enq)
			value <= value + 1'h1;
		if (reset)
			value_1 <= 1'h0;
		else if (do_deq)
			value_1 <= value_1 + 1'h1;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module TLBuffer_17 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [2:0] auto_in_a_bits_size;
	input [2:0] auto_in_a_bits_source;
	input [28:0] auto_in_a_bits_address;
	input [7:0] auto_in_a_bits_mask;
	input [63:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [2:0] auto_in_d_bits_size;
	output wire [2:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [63:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [2:0] auto_out_a_bits_size;
	output wire [2:0] auto_out_a_bits_source;
	output wire [28:0] auto_out_a_bits_address;
	output wire [7:0] auto_out_a_bits_mask;
	output wire [63:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [2:0] auto_out_d_bits_size;
	input [2:0] auto_out_d_bits_source;
	input auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [63:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [2:0] monitor_io_in_a_bits_size;
	wire [2:0] monitor_io_in_a_bits_source;
	wire [28:0] monitor_io_in_a_bits_address;
	wire [7:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_param;
	wire [2:0] monitor_io_in_d_bits_size;
	wire [2:0] monitor_io_in_d_bits_source;
	wire monitor_io_in_d_bits_sink;
	wire monitor_io_in_d_bits_denied;
	wire monitor_io_in_d_bits_corrupt;
	wire bundleOut_0_a_q_clock;
	wire bundleOut_0_a_q_reset;
	wire bundleOut_0_a_q_io_enq_ready;
	wire bundleOut_0_a_q_io_enq_valid;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_param;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_size;
	wire [2:0] bundleOut_0_a_q_io_enq_bits_source;
	wire [28:0] bundleOut_0_a_q_io_enq_bits_address;
	wire [7:0] bundleOut_0_a_q_io_enq_bits_mask;
	wire [63:0] bundleOut_0_a_q_io_enq_bits_data;
	wire bundleOut_0_a_q_io_enq_bits_corrupt;
	wire bundleOut_0_a_q_io_deq_ready;
	wire bundleOut_0_a_q_io_deq_valid;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_param;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_size;
	wire [2:0] bundleOut_0_a_q_io_deq_bits_source;
	wire [28:0] bundleOut_0_a_q_io_deq_bits_address;
	wire [7:0] bundleOut_0_a_q_io_deq_bits_mask;
	wire [63:0] bundleOut_0_a_q_io_deq_bits_data;
	wire bundleOut_0_a_q_io_deq_bits_corrupt;
	wire bundleIn_0_d_q_clock;
	wire bundleIn_0_d_q_reset;
	wire bundleIn_0_d_q_io_enq_ready;
	wire bundleIn_0_d_q_io_enq_valid;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_enq_bits_param;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_size;
	wire [2:0] bundleIn_0_d_q_io_enq_bits_source;
	wire bundleIn_0_d_q_io_enq_bits_sink;
	wire bundleIn_0_d_q_io_enq_bits_denied;
	wire [63:0] bundleIn_0_d_q_io_enq_bits_data;
	wire bundleIn_0_d_q_io_enq_bits_corrupt;
	wire bundleIn_0_d_q_io_deq_ready;
	wire bundleIn_0_d_q_io_deq_valid;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode;
	wire [1:0] bundleIn_0_d_q_io_deq_bits_param;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_size;
	wire [2:0] bundleIn_0_d_q_io_deq_bits_source;
	wire bundleIn_0_d_q_io_deq_bits_sink;
	wire bundleIn_0_d_q_io_deq_bits_denied;
	wire [63:0] bundleIn_0_d_q_io_deq_bits_data;
	wire bundleIn_0_d_q_io_deq_bits_corrupt;
	TLMonitor_45 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_param(monitor_io_in_d_bits_param),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source),
		.io_in_d_bits_sink(monitor_io_in_d_bits_sink),
		.io_in_d_bits_denied(monitor_io_in_d_bits_denied),
		.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
	);
	Queue_22 bundleOut_0_a_q(
		.clock(bundleOut_0_a_q_clock),
		.reset(bundleOut_0_a_q_reset),
		.io_enq_ready(bundleOut_0_a_q_io_enq_ready),
		.io_enq_valid(bundleOut_0_a_q_io_enq_valid),
		.io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
		.io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
		.io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
		.io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
		.io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
		.io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleOut_0_a_q_io_deq_ready),
		.io_deq_valid(bundleOut_0_a_q_io_deq_valid),
		.io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
		.io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
		.io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
		.io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
		.io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
		.io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
	);
	Queue_23 bundleIn_0_d_q(
		.clock(bundleIn_0_d_q_clock),
		.reset(bundleIn_0_d_q_reset),
		.io_enq_ready(bundleIn_0_d_q_io_enq_ready),
		.io_enq_valid(bundleIn_0_d_q_io_enq_valid),
		.io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
		.io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
		.io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
		.io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
		.io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
		.io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
		.io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
		.io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
		.io_deq_ready(bundleIn_0_d_q_io_deq_ready),
		.io_deq_valid(bundleIn_0_d_q_io_deq_valid),
		.io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
		.io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
		.io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
		.io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
		.io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
		.io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
		.io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
		.io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data;
	assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid;
	assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode;
	assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param;
	assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size;
	assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source;
	assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address;
	assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask;
	assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data;
	assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt;
	assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready;
	assign monitor_io_in_a_valid = auto_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_in_d_ready;
	assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid;
	assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode;
	assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param;
	assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size;
	assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source;
	assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink;
	assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied;
	assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt;
	assign bundleOut_0_a_q_clock = clock;
	assign bundleOut_0_a_q_reset = reset;
	assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid;
	assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode;
	assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param;
	assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size;
	assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source;
	assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address;
	assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask;
	assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data;
	assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt;
	assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready;
	assign bundleIn_0_d_q_clock = clock;
	assign bundleIn_0_d_q_reset = reset;
	assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid;
	assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode;
	assign bundleIn_0_d_q_io_enq_bits_param = auto_out_d_bits_param;
	assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size;
	assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source;
	assign bundleIn_0_d_q_io_enq_bits_sink = auto_out_d_bits_sink;
	assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied;
	assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data;
	assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt;
	assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready;
endmodule
module ClockSinkDomain_2 (
	auto_serdesser_client_out_a_ready,
	auto_serdesser_client_out_a_valid,
	auto_serdesser_client_out_a_bits_opcode,
	auto_serdesser_client_out_a_bits_param,
	auto_serdesser_client_out_a_bits_size,
	auto_serdesser_client_out_a_bits_source,
	auto_serdesser_client_out_a_bits_address,
	auto_serdesser_client_out_a_bits_mask,
	auto_serdesser_client_out_a_bits_data,
	auto_serdesser_client_out_a_bits_corrupt,
	auto_serdesser_client_out_d_ready,
	auto_serdesser_client_out_d_valid,
	auto_serdesser_client_out_d_bits_opcode,
	auto_serdesser_client_out_d_bits_param,
	auto_serdesser_client_out_d_bits_size,
	auto_serdesser_client_out_d_bits_source,
	auto_serdesser_client_out_d_bits_sink,
	auto_serdesser_client_out_d_bits_denied,
	auto_serdesser_client_out_d_bits_data,
	auto_serdesser_client_out_d_bits_corrupt,
	auto_tlserial_manager_crossing_in_a_ready,
	auto_tlserial_manager_crossing_in_a_valid,
	auto_tlserial_manager_crossing_in_a_bits_opcode,
	auto_tlserial_manager_crossing_in_a_bits_param,
	auto_tlserial_manager_crossing_in_a_bits_size,
	auto_tlserial_manager_crossing_in_a_bits_source,
	auto_tlserial_manager_crossing_in_a_bits_address,
	auto_tlserial_manager_crossing_in_a_bits_mask,
	auto_tlserial_manager_crossing_in_a_bits_data,
	auto_tlserial_manager_crossing_in_a_bits_corrupt,
	auto_tlserial_manager_crossing_in_d_ready,
	auto_tlserial_manager_crossing_in_d_valid,
	auto_tlserial_manager_crossing_in_d_bits_opcode,
	auto_tlserial_manager_crossing_in_d_bits_param,
	auto_tlserial_manager_crossing_in_d_bits_size,
	auto_tlserial_manager_crossing_in_d_bits_source,
	auto_tlserial_manager_crossing_in_d_bits_sink,
	auto_tlserial_manager_crossing_in_d_bits_denied,
	auto_tlserial_manager_crossing_in_d_bits_data,
	auto_tlserial_manager_crossing_in_d_bits_corrupt,
	auto_clock_in_clock,
	auto_clock_in_reset,
	serial_tl_in_ready,
	serial_tl_in_valid,
	serial_tl_in_bits,
	serial_tl_out_ready,
	serial_tl_out_valid,
	serial_tl_out_bits,
	clock
);
	input auto_serdesser_client_out_a_ready;
	output wire auto_serdesser_client_out_a_valid;
	output wire [2:0] auto_serdesser_client_out_a_bits_opcode;
	output wire [2:0] auto_serdesser_client_out_a_bits_param;
	output wire [3:0] auto_serdesser_client_out_a_bits_size;
	output wire auto_serdesser_client_out_a_bits_source;
	output wire [31:0] auto_serdesser_client_out_a_bits_address;
	output wire [3:0] auto_serdesser_client_out_a_bits_mask;
	output wire [31:0] auto_serdesser_client_out_a_bits_data;
	output wire auto_serdesser_client_out_a_bits_corrupt;
	output wire auto_serdesser_client_out_d_ready;
	input auto_serdesser_client_out_d_valid;
	input [2:0] auto_serdesser_client_out_d_bits_opcode;
	input [1:0] auto_serdesser_client_out_d_bits_param;
	input [3:0] auto_serdesser_client_out_d_bits_size;
	input auto_serdesser_client_out_d_bits_source;
	input auto_serdesser_client_out_d_bits_sink;
	input auto_serdesser_client_out_d_bits_denied;
	input [31:0] auto_serdesser_client_out_d_bits_data;
	input auto_serdesser_client_out_d_bits_corrupt;
	output wire auto_tlserial_manager_crossing_in_a_ready;
	input auto_tlserial_manager_crossing_in_a_valid;
	input [2:0] auto_tlserial_manager_crossing_in_a_bits_opcode;
	input [2:0] auto_tlserial_manager_crossing_in_a_bits_param;
	input [2:0] auto_tlserial_manager_crossing_in_a_bits_size;
	input [2:0] auto_tlserial_manager_crossing_in_a_bits_source;
	input [28:0] auto_tlserial_manager_crossing_in_a_bits_address;
	input [7:0] auto_tlserial_manager_crossing_in_a_bits_mask;
	input [63:0] auto_tlserial_manager_crossing_in_a_bits_data;
	input auto_tlserial_manager_crossing_in_a_bits_corrupt;
	input auto_tlserial_manager_crossing_in_d_ready;
	output wire auto_tlserial_manager_crossing_in_d_valid;
	output wire [2:0] auto_tlserial_manager_crossing_in_d_bits_opcode;
	output wire [1:0] auto_tlserial_manager_crossing_in_d_bits_param;
	output wire [2:0] auto_tlserial_manager_crossing_in_d_bits_size;
	output wire [2:0] auto_tlserial_manager_crossing_in_d_bits_source;
	output wire auto_tlserial_manager_crossing_in_d_bits_sink;
	output wire auto_tlserial_manager_crossing_in_d_bits_denied;
	output wire [63:0] auto_tlserial_manager_crossing_in_d_bits_data;
	output wire auto_tlserial_manager_crossing_in_d_bits_corrupt;
	input auto_clock_in_clock;
	input auto_clock_in_reset;
	output wire serial_tl_in_ready;
	input serial_tl_in_valid;
	input [31:0] serial_tl_in_bits;
	input serial_tl_out_ready;
	output wire serial_tl_out_valid;
	output wire [31:0] serial_tl_out_bits;
	output wire clock;
	wire serdesser_clock;
	wire serdesser_reset;
	wire serdesser_auto_manager_in_a_ready;
	wire serdesser_auto_manager_in_a_valid;
	wire [2:0] serdesser_auto_manager_in_a_bits_opcode;
	wire [2:0] serdesser_auto_manager_in_a_bits_param;
	wire [2:0] serdesser_auto_manager_in_a_bits_size;
	wire [2:0] serdesser_auto_manager_in_a_bits_source;
	wire [28:0] serdesser_auto_manager_in_a_bits_address;
	wire [7:0] serdesser_auto_manager_in_a_bits_mask;
	wire [63:0] serdesser_auto_manager_in_a_bits_data;
	wire serdesser_auto_manager_in_a_bits_corrupt;
	wire serdesser_auto_manager_in_d_ready;
	wire serdesser_auto_manager_in_d_valid;
	wire [2:0] serdesser_auto_manager_in_d_bits_opcode;
	wire [1:0] serdesser_auto_manager_in_d_bits_param;
	wire [2:0] serdesser_auto_manager_in_d_bits_size;
	wire [2:0] serdesser_auto_manager_in_d_bits_source;
	wire serdesser_auto_manager_in_d_bits_sink;
	wire serdesser_auto_manager_in_d_bits_denied;
	wire [63:0] serdesser_auto_manager_in_d_bits_data;
	wire serdesser_auto_manager_in_d_bits_corrupt;
	wire serdesser_auto_client_out_a_ready;
	wire serdesser_auto_client_out_a_valid;
	wire [2:0] serdesser_auto_client_out_a_bits_opcode;
	wire [2:0] serdesser_auto_client_out_a_bits_param;
	wire [3:0] serdesser_auto_client_out_a_bits_size;
	wire serdesser_auto_client_out_a_bits_source;
	wire [31:0] serdesser_auto_client_out_a_bits_address;
	wire [3:0] serdesser_auto_client_out_a_bits_mask;
	wire [31:0] serdesser_auto_client_out_a_bits_data;
	wire serdesser_auto_client_out_a_bits_corrupt;
	wire serdesser_auto_client_out_d_ready;
	wire serdesser_auto_client_out_d_valid;
	wire [2:0] serdesser_auto_client_out_d_bits_opcode;
	wire [1:0] serdesser_auto_client_out_d_bits_param;
	wire [3:0] serdesser_auto_client_out_d_bits_size;
	wire serdesser_auto_client_out_d_bits_source;
	wire serdesser_auto_client_out_d_bits_sink;
	wire serdesser_auto_client_out_d_bits_denied;
	wire [31:0] serdesser_auto_client_out_d_bits_data;
	wire serdesser_auto_client_out_d_bits_corrupt;
	wire serdesser_io_ser_in_ready;
	wire serdesser_io_ser_in_valid;
	wire [31:0] serdesser_io_ser_in_bits;
	wire serdesser_io_ser_out_ready;
	wire serdesser_io_ser_out_valid;
	wire [31:0] serdesser_io_ser_out_bits;
	wire buffer_clock;
	wire buffer_reset;
	wire buffer_auto_in_a_ready;
	wire buffer_auto_in_a_valid;
	wire [2:0] buffer_auto_in_a_bits_opcode;
	wire [2:0] buffer_auto_in_a_bits_param;
	wire [2:0] buffer_auto_in_a_bits_size;
	wire [2:0] buffer_auto_in_a_bits_source;
	wire [28:0] buffer_auto_in_a_bits_address;
	wire [7:0] buffer_auto_in_a_bits_mask;
	wire [63:0] buffer_auto_in_a_bits_data;
	wire buffer_auto_in_a_bits_corrupt;
	wire buffer_auto_in_d_ready;
	wire buffer_auto_in_d_valid;
	wire [2:0] buffer_auto_in_d_bits_opcode;
	wire [1:0] buffer_auto_in_d_bits_param;
	wire [2:0] buffer_auto_in_d_bits_size;
	wire [2:0] buffer_auto_in_d_bits_source;
	wire buffer_auto_in_d_bits_sink;
	wire buffer_auto_in_d_bits_denied;
	wire [63:0] buffer_auto_in_d_bits_data;
	wire buffer_auto_in_d_bits_corrupt;
	wire buffer_auto_out_a_ready;
	wire buffer_auto_out_a_valid;
	wire [2:0] buffer_auto_out_a_bits_opcode;
	wire [2:0] buffer_auto_out_a_bits_param;
	wire [2:0] buffer_auto_out_a_bits_size;
	wire [2:0] buffer_auto_out_a_bits_source;
	wire [28:0] buffer_auto_out_a_bits_address;
	wire [7:0] buffer_auto_out_a_bits_mask;
	wire [63:0] buffer_auto_out_a_bits_data;
	wire buffer_auto_out_a_bits_corrupt;
	wire buffer_auto_out_d_ready;
	wire buffer_auto_out_d_valid;
	wire [2:0] buffer_auto_out_d_bits_opcode;
	wire [1:0] buffer_auto_out_d_bits_param;
	wire [2:0] buffer_auto_out_d_bits_size;
	wire [2:0] buffer_auto_out_d_bits_source;
	wire buffer_auto_out_d_bits_sink;
	wire buffer_auto_out_d_bits_denied;
	wire [63:0] buffer_auto_out_d_bits_data;
	wire buffer_auto_out_d_bits_corrupt;
	TLSerdesser serdesser(
		.clock(serdesser_clock),
		.reset(serdesser_reset),
		.auto_manager_in_a_ready(serdesser_auto_manager_in_a_ready),
		.auto_manager_in_a_valid(serdesser_auto_manager_in_a_valid),
		.auto_manager_in_a_bits_opcode(serdesser_auto_manager_in_a_bits_opcode),
		.auto_manager_in_a_bits_param(serdesser_auto_manager_in_a_bits_param),
		.auto_manager_in_a_bits_size(serdesser_auto_manager_in_a_bits_size),
		.auto_manager_in_a_bits_source(serdesser_auto_manager_in_a_bits_source),
		.auto_manager_in_a_bits_address(serdesser_auto_manager_in_a_bits_address),
		.auto_manager_in_a_bits_mask(serdesser_auto_manager_in_a_bits_mask),
		.auto_manager_in_a_bits_data(serdesser_auto_manager_in_a_bits_data),
		.auto_manager_in_a_bits_corrupt(serdesser_auto_manager_in_a_bits_corrupt),
		.auto_manager_in_d_ready(serdesser_auto_manager_in_d_ready),
		.auto_manager_in_d_valid(serdesser_auto_manager_in_d_valid),
		.auto_manager_in_d_bits_opcode(serdesser_auto_manager_in_d_bits_opcode),
		.auto_manager_in_d_bits_param(serdesser_auto_manager_in_d_bits_param),
		.auto_manager_in_d_bits_size(serdesser_auto_manager_in_d_bits_size),
		.auto_manager_in_d_bits_source(serdesser_auto_manager_in_d_bits_source),
		.auto_manager_in_d_bits_sink(serdesser_auto_manager_in_d_bits_sink),
		.auto_manager_in_d_bits_denied(serdesser_auto_manager_in_d_bits_denied),
		.auto_manager_in_d_bits_data(serdesser_auto_manager_in_d_bits_data),
		.auto_manager_in_d_bits_corrupt(serdesser_auto_manager_in_d_bits_corrupt),
		.auto_client_out_a_ready(serdesser_auto_client_out_a_ready),
		.auto_client_out_a_valid(serdesser_auto_client_out_a_valid),
		.auto_client_out_a_bits_opcode(serdesser_auto_client_out_a_bits_opcode),
		.auto_client_out_a_bits_param(serdesser_auto_client_out_a_bits_param),
		.auto_client_out_a_bits_size(serdesser_auto_client_out_a_bits_size),
		.auto_client_out_a_bits_source(serdesser_auto_client_out_a_bits_source),
		.auto_client_out_a_bits_address(serdesser_auto_client_out_a_bits_address),
		.auto_client_out_a_bits_mask(serdesser_auto_client_out_a_bits_mask),
		.auto_client_out_a_bits_data(serdesser_auto_client_out_a_bits_data),
		.auto_client_out_a_bits_corrupt(serdesser_auto_client_out_a_bits_corrupt),
		.auto_client_out_d_ready(serdesser_auto_client_out_d_ready),
		.auto_client_out_d_valid(serdesser_auto_client_out_d_valid),
		.auto_client_out_d_bits_opcode(serdesser_auto_client_out_d_bits_opcode),
		.auto_client_out_d_bits_param(serdesser_auto_client_out_d_bits_param),
		.auto_client_out_d_bits_size(serdesser_auto_client_out_d_bits_size),
		.auto_client_out_d_bits_source(serdesser_auto_client_out_d_bits_source),
		.auto_client_out_d_bits_sink(serdesser_auto_client_out_d_bits_sink),
		.auto_client_out_d_bits_denied(serdesser_auto_client_out_d_bits_denied),
		.auto_client_out_d_bits_data(serdesser_auto_client_out_d_bits_data),
		.auto_client_out_d_bits_corrupt(serdesser_auto_client_out_d_bits_corrupt),
		.io_ser_in_ready(serdesser_io_ser_in_ready),
		.io_ser_in_valid(serdesser_io_ser_in_valid),
		.io_ser_in_bits(serdesser_io_ser_in_bits),
		.io_ser_out_ready(serdesser_io_ser_out_ready),
		.io_ser_out_valid(serdesser_io_ser_out_valid),
		.io_ser_out_bits(serdesser_io_ser_out_bits)
	);
	TLBuffer_17 buffer(
		.clock(buffer_clock),
		.reset(buffer_reset),
		.auto_in_a_ready(buffer_auto_in_a_ready),
		.auto_in_a_valid(buffer_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_auto_in_d_ready),
		.auto_in_d_valid(buffer_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(buffer_auto_in_d_bits_param),
		.auto_in_d_bits_size(buffer_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_auto_in_d_bits_source),
		.auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(buffer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(buffer_auto_out_a_ready),
		.auto_out_a_valid(buffer_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_auto_out_d_ready),
		.auto_out_d_valid(buffer_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
		.auto_out_d_bits_param(buffer_auto_out_d_bits_param),
		.auto_out_d_bits_size(buffer_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_auto_out_d_bits_source),
		.auto_out_d_bits_sink(buffer_auto_out_d_bits_sink),
		.auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
		.auto_out_d_bits_data(buffer_auto_out_d_bits_data),
		.auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt)
	);
	assign auto_serdesser_client_out_a_valid = serdesser_auto_client_out_a_valid;
	assign auto_serdesser_client_out_a_bits_opcode = serdesser_auto_client_out_a_bits_opcode;
	assign auto_serdesser_client_out_a_bits_param = serdesser_auto_client_out_a_bits_param;
	assign auto_serdesser_client_out_a_bits_size = serdesser_auto_client_out_a_bits_size;
	assign auto_serdesser_client_out_a_bits_source = serdesser_auto_client_out_a_bits_source;
	assign auto_serdesser_client_out_a_bits_address = serdesser_auto_client_out_a_bits_address;
	assign auto_serdesser_client_out_a_bits_mask = serdesser_auto_client_out_a_bits_mask;
	assign auto_serdesser_client_out_a_bits_data = serdesser_auto_client_out_a_bits_data;
	assign auto_serdesser_client_out_a_bits_corrupt = serdesser_auto_client_out_a_bits_corrupt;
	assign auto_serdesser_client_out_d_ready = serdesser_auto_client_out_d_ready;
	assign auto_tlserial_manager_crossing_in_a_ready = buffer_auto_in_a_ready;
	assign auto_tlserial_manager_crossing_in_d_valid = buffer_auto_in_d_valid;
	assign auto_tlserial_manager_crossing_in_d_bits_opcode = buffer_auto_in_d_bits_opcode;
	assign auto_tlserial_manager_crossing_in_d_bits_param = buffer_auto_in_d_bits_param;
	assign auto_tlserial_manager_crossing_in_d_bits_size = buffer_auto_in_d_bits_size;
	assign auto_tlserial_manager_crossing_in_d_bits_source = buffer_auto_in_d_bits_source;
	assign auto_tlserial_manager_crossing_in_d_bits_sink = buffer_auto_in_d_bits_sink;
	assign auto_tlserial_manager_crossing_in_d_bits_denied = buffer_auto_in_d_bits_denied;
	assign auto_tlserial_manager_crossing_in_d_bits_data = buffer_auto_in_d_bits_data;
	assign auto_tlserial_manager_crossing_in_d_bits_corrupt = buffer_auto_in_d_bits_corrupt;
	assign serial_tl_in_ready = serdesser_io_ser_in_ready;
	assign serial_tl_out_valid = serdesser_io_ser_out_valid;
	assign serial_tl_out_bits = serdesser_io_ser_out_bits;
	assign clock = auto_clock_in_clock;
	assign serdesser_clock = auto_clock_in_clock;
	assign serdesser_reset = auto_clock_in_reset;
	assign serdesser_auto_manager_in_a_valid = buffer_auto_out_a_valid;
	assign serdesser_auto_manager_in_a_bits_opcode = buffer_auto_out_a_bits_opcode;
	assign serdesser_auto_manager_in_a_bits_param = buffer_auto_out_a_bits_param;
	assign serdesser_auto_manager_in_a_bits_size = buffer_auto_out_a_bits_size;
	assign serdesser_auto_manager_in_a_bits_source = buffer_auto_out_a_bits_source;
	assign serdesser_auto_manager_in_a_bits_address = buffer_auto_out_a_bits_address;
	assign serdesser_auto_manager_in_a_bits_mask = buffer_auto_out_a_bits_mask;
	assign serdesser_auto_manager_in_a_bits_data = buffer_auto_out_a_bits_data;
	assign serdesser_auto_manager_in_a_bits_corrupt = buffer_auto_out_a_bits_corrupt;
	assign serdesser_auto_manager_in_d_ready = buffer_auto_out_d_ready;
	assign serdesser_auto_client_out_a_ready = auto_serdesser_client_out_a_ready;
	assign serdesser_auto_client_out_d_valid = auto_serdesser_client_out_d_valid;
	assign serdesser_auto_client_out_d_bits_opcode = auto_serdesser_client_out_d_bits_opcode;
	assign serdesser_auto_client_out_d_bits_param = auto_serdesser_client_out_d_bits_param;
	assign serdesser_auto_client_out_d_bits_size = auto_serdesser_client_out_d_bits_size;
	assign serdesser_auto_client_out_d_bits_source = auto_serdesser_client_out_d_bits_source;
	assign serdesser_auto_client_out_d_bits_sink = auto_serdesser_client_out_d_bits_sink;
	assign serdesser_auto_client_out_d_bits_denied = auto_serdesser_client_out_d_bits_denied;
	assign serdesser_auto_client_out_d_bits_data = auto_serdesser_client_out_d_bits_data;
	assign serdesser_auto_client_out_d_bits_corrupt = auto_serdesser_client_out_d_bits_corrupt;
	assign serdesser_io_ser_in_valid = serial_tl_in_valid;
	assign serdesser_io_ser_in_bits = serial_tl_in_bits;
	assign serdesser_io_ser_out_ready = serial_tl_out_ready;
	assign buffer_clock = auto_clock_in_clock;
	assign buffer_reset = auto_clock_in_reset;
	assign buffer_auto_in_a_valid = auto_tlserial_manager_crossing_in_a_valid;
	assign buffer_auto_in_a_bits_opcode = auto_tlserial_manager_crossing_in_a_bits_opcode;
	assign buffer_auto_in_a_bits_param = auto_tlserial_manager_crossing_in_a_bits_param;
	assign buffer_auto_in_a_bits_size = auto_tlserial_manager_crossing_in_a_bits_size;
	assign buffer_auto_in_a_bits_source = auto_tlserial_manager_crossing_in_a_bits_source;
	assign buffer_auto_in_a_bits_address = auto_tlserial_manager_crossing_in_a_bits_address;
	assign buffer_auto_in_a_bits_mask = auto_tlserial_manager_crossing_in_a_bits_mask;
	assign buffer_auto_in_a_bits_data = auto_tlserial_manager_crossing_in_a_bits_data;
	assign buffer_auto_in_a_bits_corrupt = auto_tlserial_manager_crossing_in_a_bits_corrupt;
	assign buffer_auto_in_d_ready = auto_tlserial_manager_crossing_in_d_ready;
	assign buffer_auto_out_a_ready = serdesser_auto_manager_in_a_ready;
	assign buffer_auto_out_d_valid = serdesser_auto_manager_in_d_valid;
	assign buffer_auto_out_d_bits_opcode = serdesser_auto_manager_in_d_bits_opcode;
	assign buffer_auto_out_d_bits_param = serdesser_auto_manager_in_d_bits_param;
	assign buffer_auto_out_d_bits_size = serdesser_auto_manager_in_d_bits_size;
	assign buffer_auto_out_d_bits_source = serdesser_auto_manager_in_d_bits_source;
	assign buffer_auto_out_d_bits_sink = serdesser_auto_manager_in_d_bits_sink;
	assign buffer_auto_out_d_bits_denied = serdesser_auto_manager_in_d_bits_denied;
	assign buffer_auto_out_d_bits_data = serdesser_auto_manager_in_d_bits_data;
	assign buffer_auto_out_d_bits_corrupt = serdesser_auto_manager_in_d_bits_corrupt;
endmodule
module TLBuffer_18 (
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_param,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_a_bits_corrupt,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_data,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_data
);
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [2:0] auto_in_a_bits_param;
	input [1:0] auto_in_a_bits_size;
	input [7:0] auto_in_a_bits_source;
	input [30:0] auto_in_a_bits_address;
	input [3:0] auto_in_a_bits_mask;
	input [31:0] auto_in_a_bits_data;
	input auto_in_a_bits_corrupt;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_size;
	output wire [7:0] auto_in_d_bits_source;
	output wire [31:0] auto_in_d_bits_data;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [1:0] auto_out_a_bits_size;
	output wire [7:0] auto_out_a_bits_source;
	output wire [30:0] auto_out_a_bits_address;
	output wire [3:0] auto_out_a_bits_mask;
	output wire [31:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_size;
	input [7:0] auto_out_d_bits_source;
	input [31:0] auto_out_d_bits_data;
	assign auto_in_a_ready = auto_out_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_out_a_valid = auto_in_a_valid;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_param = auto_in_a_bits_param;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module TLMonitor_46 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [1:0] io_in_a_bits_size;
	input [7:0] io_in_a_bits_source;
	input [30:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_size;
	input [7:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_4 = io_in_a_bits_source <= 8'h9f;
	wire [4:0] _is_aligned_mask_T_1 = 5'h03 << io_in_a_bits_size;
	wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0];
	wire [30:0] _GEN_71 = {29'd0, is_aligned_mask};
	wire [30:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 31'h00000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 2'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_10 = ~_source_ok_T_4;
	wire _T_20 = io_in_a_bits_opcode == 3'h6;
	wire [30:0] _T_33 = io_in_a_bits_address ^ 31'h54000000;
	wire [31:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [31:0] _T_36 = $signed(_T_34) & -32'sh00001000;
	wire _T_37 = $signed(_T_36) == 32'sh00000000;
	wire _T_69 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_73 = ~io_in_a_bits_mask;
	wire _T_74 = _T_73 == 4'h0;
	wire _T_78 = ~io_in_a_bits_corrupt;
	wire _T_82 = io_in_a_bits_opcode == 3'h7;
	wire _T_135 = io_in_a_bits_param != 3'h0;
	wire _T_148 = io_in_a_bits_opcode == 3'h4;
	wire _T_164 = io_in_a_bits_size <= 2'h2;
	wire _T_172 = _T_164 & _T_37;
	wire _T_183 = io_in_a_bits_param == 3'h0;
	wire _T_187 = io_in_a_bits_mask == mask;
	wire _T_195 = io_in_a_bits_opcode == 3'h0;
	wire _T_218 = _source_ok_T_4 & _T_172;
	wire _T_236 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_273 = ~mask;
	wire [3:0] _T_274 = io_in_a_bits_mask & _T_273;
	wire _T_275 = _T_274 == 4'h0;
	wire _T_279 = io_in_a_bits_opcode == 3'h2;
	wire _T_309 = io_in_a_bits_param <= 3'h4;
	wire _T_317 = io_in_a_bits_opcode == 3'h3;
	wire _T_347 = io_in_a_bits_param <= 3'h3;
	wire _T_355 = io_in_a_bits_opcode == 3'h5;
	wire _T_385 = io_in_a_bits_param <= 3'h1;
	wire _T_397 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_10 = io_in_d_bits_source <= 8'h9f;
	wire _T_401 = io_in_d_bits_opcode == 3'h6;
	wire _T_405 = io_in_d_bits_size >= 2'h2;
	wire _T_421 = io_in_d_bits_opcode == 3'h4;
	wire _T_449 = io_in_d_bits_opcode == 3'h5;
	wire _T_478 = io_in_d_bits_opcode == 3'h0;
	wire _T_495 = io_in_d_bits_opcode == 3'h1;
	wire _T_513 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [1:0] size;
	reg [7:0] source;
	reg [30:0] address;
	wire _T_543 = io_in_a_valid & ~a_first;
	wire _T_544 = io_in_a_bits_opcode == opcode;
	wire _T_548 = io_in_a_bits_param == param;
	wire _T_552 = io_in_a_bits_size == size;
	wire _T_556 = io_in_a_bits_source == source;
	wire _T_560 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] size_1;
	reg [7:0] source_1;
	wire _T_567 = io_in_d_valid & ~d_first;
	wire _T_568 = io_in_d_bits_opcode == opcode_1;
	wire _T_576 = io_in_d_bits_size == size_1;
	wire _T_580 = io_in_d_bits_source == source_1;
	reg [159:0] inflight;
	reg [639:0] inflight_opcodes;
	reg [639:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [10:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [639:0] _GEN_73 = {624'd0, _a_opcode_lookup_T_5};
	wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [639:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[639:1]};
	wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [639:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[639:1]};
	wire _T_594 = io_in_a_valid & a_first_1;
	wire [255:0] _a_set_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_a_bits_source;
	wire _T_597 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1;
	wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [10:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [2050:0] _GEN_1 = {2047'd0, a_opcodes_set_interm};
	wire [2050:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? _a_sizes_set_interm_T_1 : 3'h0);
	wire [2049:0] _GEN_2 = {2047'd0, a_sizes_set_interm};
	wire [2049:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [159:0] _T_599 = inflight >> io_in_a_bits_source;
	wire _T_601 = ~_T_599[0];
	wire [255:0] _GEN_16 = (a_first_done & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2050:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 2051'h0);
	wire [2049:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 2050'h0);
	wire _T_605 = io_in_d_valid & d_first_1;
	wire _T_607 = ~_T_401;
	wire _T_608 = (io_in_d_valid & d_first_1) & ~_T_401;
	wire [255:0] _d_clr_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_d_bits_source;
	wire [2062:0] _GEN_3 = {2047'd0, _a_opcode_lookup_T_5};
	wire [2062:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [255:0] _GEN_22 = ((d_first_done & d_first_1) & _T_607 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_23 = ((d_first_done & d_first_1) & _T_607 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_594 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [159:0] _T_618 = inflight >> io_in_d_bits_source;
	wire _T_620 = _T_618[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_625 = io_in_d_bits_opcode == _GEN_40;
	wire _T_626 = (io_in_d_bits_opcode == _GEN_32) | _T_625;
	wire _T_630 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_637 = io_in_d_bits_opcode == _GEN_56;
	wire _T_638 = (io_in_d_bits_opcode == _GEN_48) | _T_637;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {2'd0, io_in_d_bits_size};
	wire _T_642 = _GEN_82 == a_size_lookup;
	wire _T_652 = (((_T_605 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_607;
	wire _T_654 = ~io_in_d_ready | io_in_a_ready;
	wire [159:0] a_set = _GEN_16[159:0];
	wire [159:0] _inflight_T = inflight | a_set;
	wire [159:0] d_clr = _GEN_22[159:0];
	wire [159:0] _inflight_T_1 = ~d_clr;
	wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [639:0] a_opcodes_set = _GEN_19[639:0];
	wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [639:0] d_opcodes_clr = _GEN_23[639:0];
	wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [639:0] a_sizes_set = _GEN_20[639:0];
	wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_663 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [159:0] inflight_1;
	reg [639:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [639:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[639:1]};
	wire _T_689 = (io_in_d_valid & d_first_2) & _T_401;
	wire [255:0] _GEN_67 = ((d_first_done & d_first_2) & _T_401 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_68 = ((d_first_done & d_first_2) & _T_401 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire [159:0] _T_697 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_707 = _GEN_82 == c_size_lookup;
	wire [159:0] d_clr_1 = _GEN_67[159:0];
	wire [159:0] _inflight_T_4 = ~d_clr_1;
	wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0];
	wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_727 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			param <= io_in_a_bits_param;
		if (a_first_done & a_first)
			size <= io_in_a_bits_size;
		if (a_first_done & a_first)
			source <= io_in_a_bits_source;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 160'h0000000000000000000000000000000000000000;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 640'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 640'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 160'h0000000000000000000000000000000000000000;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 640'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (d_first_done)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module UARTTx (
	clock,
	reset,
	io_en,
	io_in_ready,
	io_in_valid,
	io_in_bits,
	io_out,
	io_div,
	io_nstop
);
	input clock;
	input reset;
	input io_en;
	output wire io_in_ready;
	input io_in_valid;
	input [7:0] io_in_bits;
	output wire io_out;
	input [15:0] io_div;
	input io_nstop;
	wire [31:0] plusarg_reader_out;
	reg [15:0] prescaler;
	wire pulse = prescaler == 16'h0000;
	reg [3:0] counter;
	reg [8:0] shifter;
	reg out;
	wire plusarg_tx = |plusarg_reader_out;
	wire busy = counter != 4'h0;
	wire _T = io_in_ready & io_in_valid;
	wire [9:0] _shifter_T_1 = {1'h1, io_in_bits, 1'h0};
	wire _counter_T = ~io_nstop;
	wire [3:0] _counter_T_2 = (_counter_T ? 4'ha : 4'h0);
	wire [3:0] _counter_T_3 = (io_nstop ? 4'hb : 4'h0);
	wire [3:0] _counter_T_4 = _counter_T_2 | _counter_T_3;
	wire [3:0] _counter_T_6 = _counter_T_4 - 4'h0;
	wire [9:0] _GEN_0 = (_T & plusarg_tx ? _shifter_T_1 : {1'd0, shifter});
	wire [15:0] _prescaler_T_2 = prescaler - 16'h0001;
	wire [3:0] _counter_T_8 = counter - 4'h1;
	wire [8:0] _shifter_T_3 = {1'h1, shifter[8:1]};
	wire [9:0] _GEN_4 = (pulse & busy ? {1'd0, _shifter_T_3} : _GEN_0);
	wire _GEN_5 = (pulse & busy ? shifter[0] : out);
	plusarg_reader #(
		.FORMAT("uart_tx=%d"),
		.DEFAULT(1),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	assign io_in_ready = io_en & ~busy;
	assign io_out = out;
	always @(posedge clock) begin
		if (reset)
			prescaler <= 16'h0000;
		else if (busy)
			if (pulse)
				prescaler <= io_div;
			else
				prescaler <= _prescaler_T_2;
		if (reset)
			counter <= 4'h0;
		else if (pulse & busy)
			counter <= _counter_T_8;
		else if (_T & plusarg_tx)
			counter <= _counter_T_6;
		shifter <= _GEN_4[8:0];
		out <= reset | _GEN_5;
	end
endmodule
module QueueCompatibility (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits,
	io_count
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [7:0] io_enq_bits;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [7:0] io_deq_bits;
	output wire [8:0] io_count;
	reg [7:0] ram [0:255];
	wire ram_io_deq_bits_MPORT_en;
	wire [7:0] ram_io_deq_bits_MPORT_addr;
	wire [7:0] ram_io_deq_bits_MPORT_data;
	wire [7:0] ram_MPORT_data;
	wire [7:0] ram_MPORT_addr;
	wire ram_MPORT_mask;
	wire ram_MPORT_en;
	reg [7:0] enq_ptr_value;
	reg [7:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = io_enq_ready & io_enq_valid;
	wire do_deq = io_deq_ready & io_deq_valid;
	wire [7:0] _value_T_1 = enq_ptr_value + 8'h01;
	wire [7:0] _value_T_3 = deq_ptr_value + 8'h01;
	wire [7:0] ptr_diff = enq_ptr_value - deq_ptr_value;
	wire [8:0] _io_count_T_1 = (maybe_full & ptr_match ? 9'h100 : 9'h000);
	wire [8:0] _GEN_11 = {1'd0, ptr_diff};
	assign ram_io_deq_bits_MPORT_en = 1'h1;
	assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
	assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr];
	assign ram_MPORT_data = io_enq_bits;
	assign ram_MPORT_addr = enq_ptr_value;
	assign ram_MPORT_mask = 1'h1;
	assign ram_MPORT_en = io_enq_ready & io_enq_valid;
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits = ram_io_deq_bits_MPORT_data;
	assign io_count = _io_count_T_1 | _GEN_11;
	always @(posedge clock) begin
		if (ram_MPORT_en & ram_MPORT_mask)
			ram[ram_MPORT_addr] <= ram_MPORT_data;
		if (reset)
			enq_ptr_value <= 8'h00;
		else if (do_enq)
			enq_ptr_value <= _value_T_1;
		if (reset)
			deq_ptr_value <= 8'h00;
		else if (do_deq)
			deq_ptr_value <= _value_T_3;
		if (reset)
			maybe_full <= 1'h0;
		else if (do_enq != do_deq)
			maybe_full <= do_enq;
	end
endmodule
module UARTRx (
	clock,
	reset,
	io_en,
	io_in,
	io_out_valid,
	io_out_bits,
	io_div
);
	input clock;
	input reset;
	input io_en;
	input io_in;
	output wire io_out_valid;
	output wire [7:0] io_out_bits;
	input [15:0] io_div;
	reg [1:0] debounce;
	wire debounce_max = debounce == 2'h3;
	wire debounce_min = debounce == 2'h0;
	reg [12:0] prescaler;
	wire pulse = prescaler == 13'h0000;
	reg [3:0] data_count;
	wire data_last = data_count == 4'h0;
	reg [3:0] sample_count;
	wire sample_mid = sample_count == 4'h7;
	wire [7:0] _countdown_T = {data_count, sample_count};
	wire [7:0] countdown = _countdown_T - 8'h01;
	wire [3:0] remainder = io_div[3:0];
	wire extend = sample_count < remainder;
	reg state;
	wire _T_5 = ~io_in;
	wire _GEN_8 = ~io_in & debounce_max;
	wire start = ~state & _GEN_8;
	wire restore = start | pulse;
	wire [12:0] prescaler_in = (restore ? {1'd0, io_div[15:4]} : prescaler);
	wire _prescaler_next_T_1 = (restore & extend ? 1'h0 : 1'h1);
	wire [12:0] _GEN_41 = {12'd0, _prescaler_next_T_1};
	wire [12:0] prescaler_next = prescaler_in - _GEN_41;
	reg [2:0] sample;
	wire _voter_T_3 = sample[0] & sample[1];
	wire _voter_T_4 = sample[0] & sample[2];
	wire _voter_T_6 = sample[1] & sample[2];
	wire voter = (_voter_T_3 | _voter_T_4) | _voter_T_6;
	reg [7:0] shifter;
	reg valid;
	wire [1:0] _debounce_T_1 = debounce - 2'h1;
	wire [1:0] _GEN_0 = (~_T_5 & ~debounce_min ? _debounce_T_1 : debounce);
	wire [1:0] _debounce_T_3 = debounce + 2'h1;
	wire [3:0] _data_count_T_3 = 4'h9 - 4'h0;
	wire _GEN_1 = debounce_max | state;
	wire [3:0] _sample_T = {sample, io_in};
	wire [7:0] _shifter_T_1 = {voter, shifter[7:1]};
	wire _GEN_12 = (data_last ? 1'h0 : state);
	wire [7:0] _GEN_14 = (data_last ? shifter : _shifter_T_1);
	wire _GEN_15 = (sample_mid ? _GEN_12 : state);
	wire _GEN_16 = sample_mid & data_last;
	wire [3:0] _GEN_18 = (pulse ? _sample_T : {1'd0, sample});
	wire _GEN_22 = pulse & _GEN_16;
	wire [3:0] _GEN_25 = (state ? _GEN_18 : {1'd0, sample});
	wire [3:0] _GEN_37 = (~state ? {1'd0, sample} : _GEN_25);
	assign io_out_valid = valid;
	assign io_out_bits = shifter;
	always @(posedge clock) begin
		if (reset)
			debounce <= 2'h0;
		else if (~io_en)
			debounce <= 2'h0;
		else if (~state)
			if (~io_in)
				debounce <= _debounce_T_3;
			else
				debounce <= _GEN_0;
		if (~state) begin
			if (~io_in)
				if (debounce_max)
					prescaler <= prescaler_next;
		end
		else if (state)
			prescaler <= prescaler_next;
		if (~state) begin
			if (~io_in)
				if (debounce_max)
					data_count <= _data_count_T_3;
		end
		else if (state)
			if (pulse)
				data_count <= countdown[7:4];
		if (~state) begin
			if (~io_in)
				if (debounce_max)
					sample_count <= 4'hf;
		end
		else if (state)
			if (pulse)
				sample_count <= countdown[3:0];
		if (reset)
			state <= 1'h0;
		else if (~state) begin
			if (~io_in)
				state <= _GEN_1;
		end
		else if (state)
			if (pulse)
				state <= _GEN_15;
		sample <= _GEN_37[2:0];
		if (!(~state))
			if (state)
				if (pulse)
					if (sample_mid)
						shifter <= _GEN_14;
		if (reset)
			valid <= 1'h0;
		else if (~state)
			valid <= 1'h0;
		else
			valid <= state & _GEN_22;
	end
endmodule
module TLUART (
	clock,
	reset,
	auto_int_xing_out_sync_0,
	auto_control_xing_in_a_ready,
	auto_control_xing_in_a_valid,
	auto_control_xing_in_a_bits_opcode,
	auto_control_xing_in_a_bits_param,
	auto_control_xing_in_a_bits_size,
	auto_control_xing_in_a_bits_source,
	auto_control_xing_in_a_bits_address,
	auto_control_xing_in_a_bits_mask,
	auto_control_xing_in_a_bits_data,
	auto_control_xing_in_a_bits_corrupt,
	auto_control_xing_in_d_ready,
	auto_control_xing_in_d_valid,
	auto_control_xing_in_d_bits_opcode,
	auto_control_xing_in_d_bits_size,
	auto_control_xing_in_d_bits_source,
	auto_control_xing_in_d_bits_data,
	auto_io_out_txd,
	auto_io_out_rxd
);
	input clock;
	input reset;
	output wire auto_int_xing_out_sync_0;
	output wire auto_control_xing_in_a_ready;
	input auto_control_xing_in_a_valid;
	input [2:0] auto_control_xing_in_a_bits_opcode;
	input [2:0] auto_control_xing_in_a_bits_param;
	input [1:0] auto_control_xing_in_a_bits_size;
	input [7:0] auto_control_xing_in_a_bits_source;
	input [30:0] auto_control_xing_in_a_bits_address;
	input [3:0] auto_control_xing_in_a_bits_mask;
	input [31:0] auto_control_xing_in_a_bits_data;
	input auto_control_xing_in_a_bits_corrupt;
	input auto_control_xing_in_d_ready;
	output wire auto_control_xing_in_d_valid;
	output wire [2:0] auto_control_xing_in_d_bits_opcode;
	output wire [1:0] auto_control_xing_in_d_bits_size;
	output wire [7:0] auto_control_xing_in_d_bits_source;
	output wire [31:0] auto_control_xing_in_d_bits_data;
	output wire auto_io_out_txd;
	input auto_io_out_rxd;
	wire buffer_auto_in_a_ready;
	wire buffer_auto_in_a_valid;
	wire [2:0] buffer_auto_in_a_bits_opcode;
	wire [2:0] buffer_auto_in_a_bits_param;
	wire [1:0] buffer_auto_in_a_bits_size;
	wire [7:0] buffer_auto_in_a_bits_source;
	wire [30:0] buffer_auto_in_a_bits_address;
	wire [3:0] buffer_auto_in_a_bits_mask;
	wire [31:0] buffer_auto_in_a_bits_data;
	wire buffer_auto_in_a_bits_corrupt;
	wire buffer_auto_in_d_ready;
	wire buffer_auto_in_d_valid;
	wire [2:0] buffer_auto_in_d_bits_opcode;
	wire [1:0] buffer_auto_in_d_bits_size;
	wire [7:0] buffer_auto_in_d_bits_source;
	wire [31:0] buffer_auto_in_d_bits_data;
	wire buffer_auto_out_a_ready;
	wire buffer_auto_out_a_valid;
	wire [2:0] buffer_auto_out_a_bits_opcode;
	wire [2:0] buffer_auto_out_a_bits_param;
	wire [1:0] buffer_auto_out_a_bits_size;
	wire [7:0] buffer_auto_out_a_bits_source;
	wire [30:0] buffer_auto_out_a_bits_address;
	wire [3:0] buffer_auto_out_a_bits_mask;
	wire [31:0] buffer_auto_out_a_bits_data;
	wire buffer_auto_out_a_bits_corrupt;
	wire buffer_auto_out_d_ready;
	wire buffer_auto_out_d_valid;
	wire [2:0] buffer_auto_out_d_bits_opcode;
	wire [1:0] buffer_auto_out_d_bits_size;
	wire [7:0] buffer_auto_out_d_bits_source;
	wire [31:0] buffer_auto_out_d_bits_data;
	wire intsource_clock;
	wire intsource_reset;
	wire intsource_auto_in_0;
	wire intsource_auto_out_sync_0;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [1:0] monitor_io_in_a_bits_size;
	wire [7:0] monitor_io_in_a_bits_source;
	wire [30:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_size;
	wire [7:0] monitor_io_in_d_bits_source;
	wire txm_clock;
	wire txm_reset;
	wire txm_io_en;
	wire txm_io_in_ready;
	wire txm_io_in_valid;
	wire [7:0] txm_io_in_bits;
	wire txm_io_out;
	wire [15:0] txm_io_div;
	wire txm_io_nstop;
	wire txq_clock;
	wire txq_reset;
	wire txq_io_enq_ready;
	wire txq_io_enq_valid;
	wire [7:0] txq_io_enq_bits;
	wire txq_io_deq_ready;
	wire txq_io_deq_valid;
	wire [7:0] txq_io_deq_bits;
	wire [8:0] txq_io_count;
	wire rxm_clock;
	wire rxm_reset;
	wire rxm_io_en;
	wire rxm_io_in;
	wire rxm_io_out_valid;
	wire [7:0] rxm_io_out_bits;
	wire [15:0] rxm_io_div;
	wire rxq_clock;
	wire rxq_reset;
	wire rxq_io_enq_ready;
	wire rxq_io_enq_valid;
	wire [7:0] rxq_io_enq_bits;
	wire rxq_io_deq_ready;
	wire rxq_io_deq_valid;
	wire [7:0] rxq_io_deq_bits;
	wire [8:0] rxq_io_count;
	reg [15:0] div;
	reg txen;
	reg rxen;
	reg [8:0] txwm;
	reg [8:0] rxwm;
	reg nstop;
	reg ie_rxwm;
	reg ie_txwm;
	wire ip_txwm = txq_io_count < txwm;
	wire ip_rxwm = rxq_io_count > rxwm;
	wire _T = ~txq_io_enq_ready;
	wire _T_1 = ~rxq_io_deq_valid;
	wire [2:0] bundleIn_0_a_bits_opcode = buffer_auto_out_a_bits_opcode;
	wire in_bits_read = bundleIn_0_a_bits_opcode == 3'h4;
	wire [30:0] bundleIn_0_a_bits_address = buffer_auto_out_a_bits_address;
	wire [9:0] in_bits_index = bundleIn_0_a_bits_address[11:2];
	wire [9:0] out_findex = in_bits_index & 10'h3f8;
	wire _out_T = out_findex == 10'h000;
	wire [3:0] bundleIn_0_a_bits_mask = buffer_auto_out_a_bits_mask;
	wire [7:0] _out_frontMask_T_5 = (bundleIn_0_a_bits_mask[0] ? 8'hff : 8'h00);
	wire [7:0] _out_frontMask_T_7 = (bundleIn_0_a_bits_mask[1] ? 8'hff : 8'h00);
	wire [7:0] _out_frontMask_T_9 = (bundleIn_0_a_bits_mask[2] ? 8'hff : 8'h00);
	wire [7:0] _out_frontMask_T_11 = (bundleIn_0_a_bits_mask[3] ? 8'hff : 8'h00);
	wire [31:0] out_frontMask = {_out_frontMask_T_11, _out_frontMask_T_9, _out_frontMask_T_7, _out_frontMask_T_5};
	wire out_rimask = |out_frontMask[7:0];
	wire out_wimask = &out_frontMask[7:0];
	wire bundleIn_0_a_valid = buffer_auto_out_a_valid;
	wire bundleIn_0_d_ready = buffer_auto_out_d_ready;
	wire [2:0] out_oindex = {in_bits_index[2], in_bits_index[1], in_bits_index[0]};
	wire [7:0] _out_frontSel_T = 8'h01 << out_oindex;
	wire out_frontSel_0 = _out_frontSel_T[0];
	wire out_wivalid_0 = (((bundleIn_0_a_valid & bundleIn_0_d_ready) & ~in_bits_read) & out_frontSel_0) & (out_findex == 10'h000);
	wire out_f_wivalid = out_wivalid_0 & out_wimask;
	wire [31:0] bundleIn_0_a_bits_data = buffer_auto_out_a_bits_data;
	wire out_womask_2 = &out_frontMask[31];
	wire out_f_woready_2 = out_wivalid_0 & out_womask_2;
	wire quash = out_f_woready_2 & bundleIn_0_a_bits_data[31];
	wire [31:0] out_prepend_1 = {_T, 31'h00000000};
	wire out_wimask_3 = &out_frontMask[0];
	wire out_wimask_4 = &out_frontMask[1];
	wire [1:0] out_prepend_2 = {ip_rxwm, ip_txwm};
	wire out_frontSel_1 = _out_frontSel_T[1];
	wire out_rivalid_5 = (((bundleIn_0_a_valid & bundleIn_0_d_ready) & in_bits_read) & out_frontSel_1) & (out_findex == 10'h000);
	wire [7:0] _out_T_66 = rxq_io_deq_bits;
	wire [8:0] out_prepend_3 = {1'h0, _out_T_66};
	wire [30:0] _out_T_75 = {22'd0, out_prepend_3};
	wire [31:0] out_prepend_4 = {_T_1, _out_T_75};
	wire out_wimask_8 = &out_frontMask[15:0];
	wire out_frontSel_6 = _out_frontSel_T[6];
	wire out_wivalid_8 = (((bundleIn_0_a_valid & bundleIn_0_d_ready) & ~in_bits_read) & out_frontSel_6) & (out_findex == 10'h000);
	wire out_f_wivalid_8 = out_wivalid_8 & out_wimask_8;
	wire out_frontSel_2 = _out_frontSel_T[2];
	wire out_wivalid_9 = (((bundleIn_0_a_valid & bundleIn_0_d_ready) & ~in_bits_read) & out_frontSel_2) & (out_findex == 10'h000);
	wire out_f_wivalid_9 = out_wivalid_9 & out_wimask_3;
	wire out_f_wivalid_10 = out_wivalid_9 & out_wimask_4;
	wire [1:0] out_prepend_5 = {nstop, txen};
	wire out_wimask_11 = &out_frontMask[24:16];
	wire out_f_wivalid_11 = out_wivalid_9 & out_wimask_11;
	wire [15:0] _out_prepend_T_6 = {14'd0, out_prepend_5};
	wire [24:0] out_prepend_6 = {txwm, _out_prepend_T_6};
	wire out_frontSel_3 = _out_frontSel_T[3];
	wire out_wivalid_12 = (((bundleIn_0_a_valid & bundleIn_0_d_ready) & ~in_bits_read) & out_frontSel_3) & (out_findex == 10'h000);
	wire out_f_wivalid_12 = out_wivalid_12 & out_wimask_3;
	wire out_f_wivalid_13 = out_wivalid_12 & out_wimask_11;
	wire [15:0] _out_prepend_T_7 = {15'd0, rxen};
	wire [24:0] out_prepend_7 = {rxwm, _out_prepend_T_7};
	wire out_frontSel_4 = _out_frontSel_T[4];
	wire out_wivalid_14 = (((bundleIn_0_a_valid & bundleIn_0_d_ready) & ~in_bits_read) & out_frontSel_4) & (out_findex == 10'h000);
	wire out_f_wivalid_14 = out_wivalid_14 & out_wimask_3;
	wire out_f_wivalid_15 = out_wivalid_14 & out_wimask_4;
	wire [1:0] out_prepend_8 = {ie_rxwm, ie_txwm};
	wire _GEN_41 = (3'h1 == out_oindex ? _out_T : _out_T);
	wire _GEN_42 = (3'h2 == out_oindex ? _out_T : _GEN_41);
	wire _GEN_43 = (3'h3 == out_oindex ? _out_T : _GEN_42);
	wire _GEN_44 = (3'h4 == out_oindex ? _out_T : _GEN_43);
	wire _GEN_45 = (3'h5 == out_oindex ? _out_T : _GEN_44);
	wire _GEN_46 = (3'h6 == out_oindex ? _out_T : _GEN_45);
	wire _GEN_47 = (3'h7 == out_oindex) | _GEN_46;
	wire [31:0] _GEN_49 = (3'h1 == out_oindex ? out_prepend_4 : out_prepend_1);
	wire [31:0] _out_out_bits_data_WIRE_1_2 = {7'd0, out_prepend_6};
	wire [31:0] _GEN_50 = (3'h2 == out_oindex ? _out_out_bits_data_WIRE_1_2 : _GEN_49);
	wire [31:0] _out_out_bits_data_WIRE_1_3 = {7'd0, out_prepend_7};
	wire [31:0] _GEN_51 = (3'h3 == out_oindex ? _out_out_bits_data_WIRE_1_3 : _GEN_50);
	wire [31:0] _out_out_bits_data_WIRE_1_4 = {30'd0, out_prepend_8};
	wire [31:0] _GEN_52 = (3'h4 == out_oindex ? _out_out_bits_data_WIRE_1_4 : _GEN_51);
	wire [31:0] _out_out_bits_data_WIRE_1_5 = {30'd0, out_prepend_2};
	wire [31:0] _GEN_53 = (3'h5 == out_oindex ? _out_out_bits_data_WIRE_1_5 : _GEN_52);
	wire [31:0] _out_out_bits_data_WIRE_1_6 = {16'd0, div};
	wire [31:0] _GEN_54 = (3'h6 == out_oindex ? _out_out_bits_data_WIRE_1_6 : _GEN_53);
	wire [31:0] _GEN_55 = (3'h7 == out_oindex ? 32'h00000000 : _GEN_54);
	TLBuffer_18 buffer(
		.auto_in_a_ready(buffer_auto_in_a_ready),
		.auto_in_a_valid(buffer_auto_in_a_valid),
		.auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(buffer_auto_in_a_bits_param),
		.auto_in_a_bits_size(buffer_auto_in_a_bits_size),
		.auto_in_a_bits_source(buffer_auto_in_a_bits_source),
		.auto_in_a_bits_address(buffer_auto_in_a_bits_address),
		.auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
		.auto_in_a_bits_data(buffer_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
		.auto_in_d_ready(buffer_auto_in_d_ready),
		.auto_in_d_valid(buffer_auto_in_d_valid),
		.auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(buffer_auto_in_d_bits_size),
		.auto_in_d_bits_source(buffer_auto_in_d_bits_source),
		.auto_in_d_bits_data(buffer_auto_in_d_bits_data),
		.auto_out_a_ready(buffer_auto_out_a_ready),
		.auto_out_a_valid(buffer_auto_out_a_valid),
		.auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
		.auto_out_a_bits_param(buffer_auto_out_a_bits_param),
		.auto_out_a_bits_size(buffer_auto_out_a_bits_size),
		.auto_out_a_bits_source(buffer_auto_out_a_bits_source),
		.auto_out_a_bits_address(buffer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(buffer_auto_out_a_bits_data),
		.auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
		.auto_out_d_ready(buffer_auto_out_d_ready),
		.auto_out_d_valid(buffer_auto_out_d_valid),
		.auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
		.auto_out_d_bits_size(buffer_auto_out_d_bits_size),
		.auto_out_d_bits_source(buffer_auto_out_d_bits_source),
		.auto_out_d_bits_data(buffer_auto_out_d_bits_data)
	);
	IntSyncCrossingSource_1 intsource(
		.clock(intsource_clock),
		.reset(intsource_reset),
		.auto_in_0(intsource_auto_in_0),
		.auto_out_sync_0(intsource_auto_out_sync_0)
	);
	TLMonitor_46 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	UARTTx txm(
		.clock(txm_clock),
		.reset(txm_reset),
		.io_en(txm_io_en),
		.io_in_ready(txm_io_in_ready),
		.io_in_valid(txm_io_in_valid),
		.io_in_bits(txm_io_in_bits),
		.io_out(txm_io_out),
		.io_div(txm_io_div),
		.io_nstop(txm_io_nstop)
	);
	QueueCompatibility txq(
		.clock(txq_clock),
		.reset(txq_reset),
		.io_enq_ready(txq_io_enq_ready),
		.io_enq_valid(txq_io_enq_valid),
		.io_enq_bits(txq_io_enq_bits),
		.io_deq_ready(txq_io_deq_ready),
		.io_deq_valid(txq_io_deq_valid),
		.io_deq_bits(txq_io_deq_bits),
		.io_count(txq_io_count)
	);
	UARTRx rxm(
		.clock(rxm_clock),
		.reset(rxm_reset),
		.io_en(rxm_io_en),
		.io_in(rxm_io_in),
		.io_out_valid(rxm_io_out_valid),
		.io_out_bits(rxm_io_out_bits),
		.io_div(rxm_io_div)
	);
	QueueCompatibility rxq(
		.clock(rxq_clock),
		.reset(rxq_reset),
		.io_enq_ready(rxq_io_enq_ready),
		.io_enq_valid(rxq_io_enq_valid),
		.io_enq_bits(rxq_io_enq_bits),
		.io_deq_ready(rxq_io_deq_ready),
		.io_deq_valid(rxq_io_deq_valid),
		.io_deq_bits(rxq_io_deq_bits),
		.io_count(rxq_io_count)
	);
	assign auto_int_xing_out_sync_0 = intsource_auto_out_sync_0;
	assign auto_control_xing_in_a_ready = buffer_auto_in_a_ready;
	assign auto_control_xing_in_d_valid = buffer_auto_in_d_valid;
	assign auto_control_xing_in_d_bits_opcode = buffer_auto_in_d_bits_opcode;
	assign auto_control_xing_in_d_bits_size = buffer_auto_in_d_bits_size;
	assign auto_control_xing_in_d_bits_source = buffer_auto_in_d_bits_source;
	assign auto_control_xing_in_d_bits_data = buffer_auto_in_d_bits_data;
	assign auto_io_out_txd = txm_io_out;
	assign buffer_auto_in_a_valid = auto_control_xing_in_a_valid;
	assign buffer_auto_in_a_bits_opcode = auto_control_xing_in_a_bits_opcode;
	assign buffer_auto_in_a_bits_param = auto_control_xing_in_a_bits_param;
	assign buffer_auto_in_a_bits_size = auto_control_xing_in_a_bits_size;
	assign buffer_auto_in_a_bits_source = auto_control_xing_in_a_bits_source;
	assign buffer_auto_in_a_bits_address = auto_control_xing_in_a_bits_address;
	assign buffer_auto_in_a_bits_mask = auto_control_xing_in_a_bits_mask;
	assign buffer_auto_in_a_bits_data = auto_control_xing_in_a_bits_data;
	assign buffer_auto_in_a_bits_corrupt = auto_control_xing_in_a_bits_corrupt;
	assign buffer_auto_in_d_ready = auto_control_xing_in_d_ready;
	assign buffer_auto_out_a_ready = buffer_auto_out_d_ready;
	assign buffer_auto_out_d_valid = buffer_auto_out_a_valid;
	assign buffer_auto_out_d_bits_opcode = {2'd0, in_bits_read};
	assign buffer_auto_out_d_bits_size = buffer_auto_out_a_bits_size;
	assign buffer_auto_out_d_bits_source = buffer_auto_out_a_bits_source;
	assign buffer_auto_out_d_bits_data = (_GEN_47 ? _GEN_55 : 32'h00000000);
	assign intsource_clock = clock;
	assign intsource_reset = reset;
	assign intsource_auto_in_0 = (ip_txwm & ie_txwm) | (ip_rxwm & ie_rxwm);
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = buffer_auto_out_d_ready;
	assign monitor_io_in_a_valid = buffer_auto_out_a_valid;
	assign monitor_io_in_a_bits_opcode = buffer_auto_out_a_bits_opcode;
	assign monitor_io_in_a_bits_param = buffer_auto_out_a_bits_param;
	assign monitor_io_in_a_bits_size = buffer_auto_out_a_bits_size;
	assign monitor_io_in_a_bits_source = buffer_auto_out_a_bits_source;
	assign monitor_io_in_a_bits_address = buffer_auto_out_a_bits_address;
	assign monitor_io_in_a_bits_mask = buffer_auto_out_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = buffer_auto_out_a_bits_corrupt;
	assign monitor_io_in_d_ready = buffer_auto_out_d_ready;
	assign monitor_io_in_d_valid = buffer_auto_out_a_valid;
	assign monitor_io_in_d_bits_opcode = {2'd0, in_bits_read};
	assign monitor_io_in_d_bits_size = buffer_auto_out_a_bits_size;
	assign monitor_io_in_d_bits_source = buffer_auto_out_a_bits_source;
	assign txm_clock = clock;
	assign txm_reset = reset;
	assign txm_io_en = txen;
	assign txm_io_in_valid = txq_io_deq_valid;
	assign txm_io_in_bits = txq_io_deq_bits;
	assign txm_io_div = div;
	assign txm_io_nstop = nstop;
	assign txq_clock = clock;
	assign txq_reset = reset;
	assign txq_io_enq_valid = out_f_wivalid & ~quash;
	assign txq_io_enq_bits = bundleIn_0_a_bits_data[7:0];
	assign txq_io_deq_ready = txm_io_in_ready;
	assign rxm_clock = clock;
	assign rxm_reset = reset;
	assign rxm_io_en = rxen;
	assign rxm_io_in = auto_io_out_rxd;
	assign rxm_io_div = div;
	assign rxq_clock = clock;
	assign rxq_reset = reset;
	assign rxq_io_enq_valid = rxm_io_out_valid;
	assign rxq_io_enq_bits = rxm_io_out_bits;
	assign rxq_io_deq_ready = out_rivalid_5 & out_rimask;
	always @(posedge clock) begin
		if (reset)
			div <= 16'h0364;
		else if (out_f_wivalid_8)
			div <= bundleIn_0_a_bits_data[15:0];
		if (reset)
			txen <= 1'h0;
		else if (out_f_wivalid_9)
			txen <= bundleIn_0_a_bits_data[0];
		if (reset)
			rxen <= 1'h0;
		else if (out_f_wivalid_12)
			rxen <= bundleIn_0_a_bits_data[0];
		if (reset)
			txwm <= 9'h000;
		else if (out_f_wivalid_11)
			txwm <= bundleIn_0_a_bits_data[24:16];
		if (reset)
			rxwm <= 9'h000;
		else if (out_f_wivalid_13)
			rxwm <= bundleIn_0_a_bits_data[24:16];
		if (reset)
			nstop <= 1'h0;
		else if (out_f_wivalid_10)
			nstop <= bundleIn_0_a_bits_data[1];
		if (reset)
			ie_rxwm <= 1'h0;
		else if (out_f_wivalid_15)
			ie_rxwm <= bundleIn_0_a_bits_data[1];
		if (reset)
			ie_txwm <= 1'h0;
		else if (out_f_wivalid_14)
			ie_txwm <= bundleIn_0_a_bits_data[0];
	end
endmodule
module ClockSinkDomain_3 (
	auto_uart_0_int_xing_out_sync_0,
	auto_uart_0_control_xing_in_a_ready,
	auto_uart_0_control_xing_in_a_valid,
	auto_uart_0_control_xing_in_a_bits_opcode,
	auto_uart_0_control_xing_in_a_bits_param,
	auto_uart_0_control_xing_in_a_bits_size,
	auto_uart_0_control_xing_in_a_bits_source,
	auto_uart_0_control_xing_in_a_bits_address,
	auto_uart_0_control_xing_in_a_bits_mask,
	auto_uart_0_control_xing_in_a_bits_data,
	auto_uart_0_control_xing_in_a_bits_corrupt,
	auto_uart_0_control_xing_in_d_ready,
	auto_uart_0_control_xing_in_d_valid,
	auto_uart_0_control_xing_in_d_bits_opcode,
	auto_uart_0_control_xing_in_d_bits_size,
	auto_uart_0_control_xing_in_d_bits_source,
	auto_uart_0_control_xing_in_d_bits_data,
	auto_uart_0_io_out_txd,
	auto_uart_0_io_out_rxd,
	auto_clock_in_clock,
	auto_clock_in_reset
);
	output wire auto_uart_0_int_xing_out_sync_0;
	output wire auto_uart_0_control_xing_in_a_ready;
	input auto_uart_0_control_xing_in_a_valid;
	input [2:0] auto_uart_0_control_xing_in_a_bits_opcode;
	input [2:0] auto_uart_0_control_xing_in_a_bits_param;
	input [1:0] auto_uart_0_control_xing_in_a_bits_size;
	input [7:0] auto_uart_0_control_xing_in_a_bits_source;
	input [30:0] auto_uart_0_control_xing_in_a_bits_address;
	input [3:0] auto_uart_0_control_xing_in_a_bits_mask;
	input [31:0] auto_uart_0_control_xing_in_a_bits_data;
	input auto_uart_0_control_xing_in_a_bits_corrupt;
	input auto_uart_0_control_xing_in_d_ready;
	output wire auto_uart_0_control_xing_in_d_valid;
	output wire [2:0] auto_uart_0_control_xing_in_d_bits_opcode;
	output wire [1:0] auto_uart_0_control_xing_in_d_bits_size;
	output wire [7:0] auto_uart_0_control_xing_in_d_bits_source;
	output wire [31:0] auto_uart_0_control_xing_in_d_bits_data;
	output wire auto_uart_0_io_out_txd;
	input auto_uart_0_io_out_rxd;
	input auto_clock_in_clock;
	input auto_clock_in_reset;
	wire uart_0_clock;
	wire uart_0_reset;
	wire uart_0_auto_int_xing_out_sync_0;
	wire uart_0_auto_control_xing_in_a_ready;
	wire uart_0_auto_control_xing_in_a_valid;
	wire [2:0] uart_0_auto_control_xing_in_a_bits_opcode;
	wire [2:0] uart_0_auto_control_xing_in_a_bits_param;
	wire [1:0] uart_0_auto_control_xing_in_a_bits_size;
	wire [7:0] uart_0_auto_control_xing_in_a_bits_source;
	wire [30:0] uart_0_auto_control_xing_in_a_bits_address;
	wire [3:0] uart_0_auto_control_xing_in_a_bits_mask;
	wire [31:0] uart_0_auto_control_xing_in_a_bits_data;
	wire uart_0_auto_control_xing_in_a_bits_corrupt;
	wire uart_0_auto_control_xing_in_d_ready;
	wire uart_0_auto_control_xing_in_d_valid;
	wire [2:0] uart_0_auto_control_xing_in_d_bits_opcode;
	wire [1:0] uart_0_auto_control_xing_in_d_bits_size;
	wire [7:0] uart_0_auto_control_xing_in_d_bits_source;
	wire [31:0] uart_0_auto_control_xing_in_d_bits_data;
	wire uart_0_auto_io_out_txd;
	wire uart_0_auto_io_out_rxd;
	TLUART uart_0(
		.clock(uart_0_clock),
		.reset(uart_0_reset),
		.auto_int_xing_out_sync_0(uart_0_auto_int_xing_out_sync_0),
		.auto_control_xing_in_a_ready(uart_0_auto_control_xing_in_a_ready),
		.auto_control_xing_in_a_valid(uart_0_auto_control_xing_in_a_valid),
		.auto_control_xing_in_a_bits_opcode(uart_0_auto_control_xing_in_a_bits_opcode),
		.auto_control_xing_in_a_bits_param(uart_0_auto_control_xing_in_a_bits_param),
		.auto_control_xing_in_a_bits_size(uart_0_auto_control_xing_in_a_bits_size),
		.auto_control_xing_in_a_bits_source(uart_0_auto_control_xing_in_a_bits_source),
		.auto_control_xing_in_a_bits_address(uart_0_auto_control_xing_in_a_bits_address),
		.auto_control_xing_in_a_bits_mask(uart_0_auto_control_xing_in_a_bits_mask),
		.auto_control_xing_in_a_bits_data(uart_0_auto_control_xing_in_a_bits_data),
		.auto_control_xing_in_a_bits_corrupt(uart_0_auto_control_xing_in_a_bits_corrupt),
		.auto_control_xing_in_d_ready(uart_0_auto_control_xing_in_d_ready),
		.auto_control_xing_in_d_valid(uart_0_auto_control_xing_in_d_valid),
		.auto_control_xing_in_d_bits_opcode(uart_0_auto_control_xing_in_d_bits_opcode),
		.auto_control_xing_in_d_bits_size(uart_0_auto_control_xing_in_d_bits_size),
		.auto_control_xing_in_d_bits_source(uart_0_auto_control_xing_in_d_bits_source),
		.auto_control_xing_in_d_bits_data(uart_0_auto_control_xing_in_d_bits_data),
		.auto_io_out_txd(uart_0_auto_io_out_txd),
		.auto_io_out_rxd(uart_0_auto_io_out_rxd)
	);
	assign auto_uart_0_int_xing_out_sync_0 = uart_0_auto_int_xing_out_sync_0;
	assign auto_uart_0_control_xing_in_a_ready = uart_0_auto_control_xing_in_a_ready;
	assign auto_uart_0_control_xing_in_d_valid = uart_0_auto_control_xing_in_d_valid;
	assign auto_uart_0_control_xing_in_d_bits_opcode = uart_0_auto_control_xing_in_d_bits_opcode;
	assign auto_uart_0_control_xing_in_d_bits_size = uart_0_auto_control_xing_in_d_bits_size;
	assign auto_uart_0_control_xing_in_d_bits_source = uart_0_auto_control_xing_in_d_bits_source;
	assign auto_uart_0_control_xing_in_d_bits_data = uart_0_auto_control_xing_in_d_bits_data;
	assign auto_uart_0_io_out_txd = uart_0_auto_io_out_txd;
	assign uart_0_clock = auto_clock_in_clock;
	assign uart_0_reset = auto_clock_in_reset;
	assign uart_0_auto_control_xing_in_a_valid = auto_uart_0_control_xing_in_a_valid;
	assign uart_0_auto_control_xing_in_a_bits_opcode = auto_uart_0_control_xing_in_a_bits_opcode;
	assign uart_0_auto_control_xing_in_a_bits_param = auto_uart_0_control_xing_in_a_bits_param;
	assign uart_0_auto_control_xing_in_a_bits_size = auto_uart_0_control_xing_in_a_bits_size;
	assign uart_0_auto_control_xing_in_a_bits_source = auto_uart_0_control_xing_in_a_bits_source;
	assign uart_0_auto_control_xing_in_a_bits_address = auto_uart_0_control_xing_in_a_bits_address;
	assign uart_0_auto_control_xing_in_a_bits_mask = auto_uart_0_control_xing_in_a_bits_mask;
	assign uart_0_auto_control_xing_in_a_bits_data = auto_uart_0_control_xing_in_a_bits_data;
	assign uart_0_auto_control_xing_in_a_bits_corrupt = auto_uart_0_control_xing_in_a_bits_corrupt;
	assign uart_0_auto_control_xing_in_d_ready = auto_uart_0_control_xing_in_d_ready;
	assign uart_0_auto_io_out_rxd = auto_uart_0_io_out_rxd;
endmodule
module TLMonitor_47 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [1:0] io_in_a_bits_size;
	input [7:0] io_in_a_bits_source;
	input [20:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_size;
	input [7:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_4 = io_in_a_bits_source <= 8'h9f;
	wire [4:0] _is_aligned_mask_T_1 = 5'h03 << io_in_a_bits_size;
	wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0];
	wire [20:0] _GEN_71 = {19'd0, is_aligned_mask};
	wire [20:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 21'h000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 2'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_10 = ~_source_ok_T_4;
	wire _T_20 = io_in_a_bits_opcode == 3'h6;
	wire [20:0] _T_33 = io_in_a_bits_address ^ 21'h100000;
	wire [21:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [21:0] _T_36 = $signed(_T_34) & -22'sh001000;
	wire _T_37 = $signed(_T_36) == 22'sh000000;
	wire _T_69 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_73 = ~io_in_a_bits_mask;
	wire _T_74 = _T_73 == 4'h0;
	wire _T_78 = ~io_in_a_bits_corrupt;
	wire _T_82 = io_in_a_bits_opcode == 3'h7;
	wire _T_135 = io_in_a_bits_param != 3'h0;
	wire _T_148 = io_in_a_bits_opcode == 3'h4;
	wire _T_164 = io_in_a_bits_size <= 2'h2;
	wire _T_172 = _T_164 & _T_37;
	wire _T_183 = io_in_a_bits_param == 3'h0;
	wire _T_187 = io_in_a_bits_mask == mask;
	wire _T_195 = io_in_a_bits_opcode == 3'h0;
	wire _T_218 = _source_ok_T_4 & _T_172;
	wire _T_236 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_273 = ~mask;
	wire [3:0] _T_274 = io_in_a_bits_mask & _T_273;
	wire _T_275 = _T_274 == 4'h0;
	wire _T_279 = io_in_a_bits_opcode == 3'h2;
	wire _T_309 = io_in_a_bits_param <= 3'h4;
	wire _T_317 = io_in_a_bits_opcode == 3'h3;
	wire _T_347 = io_in_a_bits_param <= 3'h3;
	wire _T_355 = io_in_a_bits_opcode == 3'h5;
	wire _T_385 = io_in_a_bits_param <= 3'h1;
	wire _T_397 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_10 = io_in_d_bits_source <= 8'h9f;
	wire _T_401 = io_in_d_bits_opcode == 3'h6;
	wire _T_405 = io_in_d_bits_size >= 2'h2;
	wire _T_421 = io_in_d_bits_opcode == 3'h4;
	wire _T_449 = io_in_d_bits_opcode == 3'h5;
	wire _T_478 = io_in_d_bits_opcode == 3'h0;
	wire _T_495 = io_in_d_bits_opcode == 3'h1;
	wire _T_513 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [1:0] size;
	reg [7:0] source;
	reg [20:0] address;
	wire _T_543 = io_in_a_valid & ~a_first;
	wire _T_544 = io_in_a_bits_opcode == opcode;
	wire _T_548 = io_in_a_bits_param == param;
	wire _T_552 = io_in_a_bits_size == size;
	wire _T_556 = io_in_a_bits_source == source;
	wire _T_560 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] size_1;
	reg [7:0] source_1;
	wire _T_567 = io_in_d_valid & ~d_first;
	wire _T_568 = io_in_d_bits_opcode == opcode_1;
	wire _T_576 = io_in_d_bits_size == size_1;
	wire _T_580 = io_in_d_bits_source == source_1;
	reg [159:0] inflight;
	reg [639:0] inflight_opcodes;
	reg [639:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [10:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [639:0] _GEN_73 = {624'd0, _a_opcode_lookup_T_5};
	wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [639:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[639:1]};
	wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [639:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[639:1]};
	wire _T_594 = io_in_a_valid & a_first_1;
	wire [255:0] _a_set_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_a_bits_source;
	wire _T_597 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1;
	wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [10:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [2050:0] _GEN_1 = {2047'd0, a_opcodes_set_interm};
	wire [2050:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? _a_sizes_set_interm_T_1 : 3'h0);
	wire [2049:0] _GEN_2 = {2047'd0, a_sizes_set_interm};
	wire [2049:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [159:0] _T_599 = inflight >> io_in_a_bits_source;
	wire _T_601 = ~_T_599[0];
	wire [255:0] _GEN_16 = (a_first_done & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2050:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 2051'h0);
	wire [2049:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 2050'h0);
	wire _T_605 = io_in_d_valid & d_first_1;
	wire _T_607 = ~_T_401;
	wire _T_608 = (io_in_d_valid & d_first_1) & ~_T_401;
	wire [255:0] _d_clr_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_d_bits_source;
	wire [2062:0] _GEN_3 = {2047'd0, _a_opcode_lookup_T_5};
	wire [2062:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [255:0] _GEN_22 = ((d_first_done & d_first_1) & _T_607 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_23 = ((d_first_done & d_first_1) & _T_607 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_594 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [159:0] _T_618 = inflight >> io_in_d_bits_source;
	wire _T_620 = _T_618[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_625 = io_in_d_bits_opcode == _GEN_40;
	wire _T_626 = (io_in_d_bits_opcode == _GEN_32) | _T_625;
	wire _T_630 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_637 = io_in_d_bits_opcode == _GEN_56;
	wire _T_638 = (io_in_d_bits_opcode == _GEN_48) | _T_637;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {2'd0, io_in_d_bits_size};
	wire _T_642 = _GEN_82 == a_size_lookup;
	wire _T_652 = (((_T_605 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_607;
	wire _T_654 = ~io_in_d_ready | io_in_a_ready;
	wire [159:0] a_set = _GEN_16[159:0];
	wire [159:0] _inflight_T = inflight | a_set;
	wire [159:0] d_clr = _GEN_22[159:0];
	wire [159:0] _inflight_T_1 = ~d_clr;
	wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [639:0] a_opcodes_set = _GEN_19[639:0];
	wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [639:0] d_opcodes_clr = _GEN_23[639:0];
	wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [639:0] a_sizes_set = _GEN_20[639:0];
	wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_663 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [159:0] inflight_1;
	reg [639:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [639:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[639:1]};
	wire _T_689 = (io_in_d_valid & d_first_2) & _T_401;
	wire [255:0] _GEN_67 = ((d_first_done & d_first_2) & _T_401 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_68 = ((d_first_done & d_first_2) & _T_401 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire [159:0] _T_697 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_707 = _GEN_82 == c_size_lookup;
	wire [159:0] d_clr_1 = _GEN_67[159:0];
	wire [159:0] _inflight_T_4 = ~d_clr_1;
	wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0];
	wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_727 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			param <= io_in_a_bits_param;
		if (a_first_done & a_first)
			size <= io_in_a_bits_size;
		if (a_first_done & a_first)
			source <= io_in_a_bits_source;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 160'h0000000000000000000000000000000000000000;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 640'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 640'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 160'h0000000000000000000000000000000000000000;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 640'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (d_first_done)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module AsyncResetRegVec_w1_i1 (
	clock,
	reset,
	io_d,
	io_q,
	io_en
);
	input clock;
	input reset;
	input io_d;
	output wire io_q;
	input io_en;
	reg reg_;
	assign io_q = reg_;
	always @(posedge clock or posedge reset)
		if (reset)
			reg_ <= 1'h1;
		else if (io_en)
			reg_ <= io_d;
endmodule
module TileClockGater (
	clock,
	reset,
	auto_tile_clock_gater_in_1_a_ready,
	auto_tile_clock_gater_in_1_a_valid,
	auto_tile_clock_gater_in_1_a_bits_opcode,
	auto_tile_clock_gater_in_1_a_bits_param,
	auto_tile_clock_gater_in_1_a_bits_size,
	auto_tile_clock_gater_in_1_a_bits_source,
	auto_tile_clock_gater_in_1_a_bits_address,
	auto_tile_clock_gater_in_1_a_bits_mask,
	auto_tile_clock_gater_in_1_a_bits_data,
	auto_tile_clock_gater_in_1_a_bits_corrupt,
	auto_tile_clock_gater_in_1_d_ready,
	auto_tile_clock_gater_in_1_d_valid,
	auto_tile_clock_gater_in_1_d_bits_opcode,
	auto_tile_clock_gater_in_1_d_bits_size,
	auto_tile_clock_gater_in_1_d_bits_source,
	auto_tile_clock_gater_in_1_d_bits_data,
	auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_clock,
	auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_reset,
	auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_clock,
	auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_reset,
	auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_clock,
	auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_reset,
	auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_clock,
	auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_reset,
	auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_clock,
	auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_reset,
	auto_tile_clock_gater_out_member_allClocks_implicit_clock_clock,
	auto_tile_clock_gater_out_member_allClocks_implicit_clock_reset,
	auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock,
	auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset,
	auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock,
	auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset,
	auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock,
	auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset,
	auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock,
	auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset
);
	input clock;
	input reset;
	output wire auto_tile_clock_gater_in_1_a_ready;
	input auto_tile_clock_gater_in_1_a_valid;
	input [2:0] auto_tile_clock_gater_in_1_a_bits_opcode;
	input [2:0] auto_tile_clock_gater_in_1_a_bits_param;
	input [1:0] auto_tile_clock_gater_in_1_a_bits_size;
	input [7:0] auto_tile_clock_gater_in_1_a_bits_source;
	input [20:0] auto_tile_clock_gater_in_1_a_bits_address;
	input [3:0] auto_tile_clock_gater_in_1_a_bits_mask;
	input [31:0] auto_tile_clock_gater_in_1_a_bits_data;
	input auto_tile_clock_gater_in_1_a_bits_corrupt;
	input auto_tile_clock_gater_in_1_d_ready;
	output wire auto_tile_clock_gater_in_1_d_valid;
	output wire [2:0] auto_tile_clock_gater_in_1_d_bits_opcode;
	output wire [1:0] auto_tile_clock_gater_in_1_d_bits_size;
	output wire [7:0] auto_tile_clock_gater_in_1_d_bits_source;
	output wire [31:0] auto_tile_clock_gater_in_1_d_bits_data;
	input auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_clock;
	input auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_reset;
	input auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_clock;
	input auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_reset;
	input auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_clock;
	input auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_reset;
	input auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_clock;
	input auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_reset;
	input auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_clock;
	input auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_reset;
	output wire auto_tile_clock_gater_out_member_allClocks_implicit_clock_clock;
	output wire auto_tile_clock_gater_out_member_allClocks_implicit_clock_reset;
	output wire auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock;
	output wire auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset;
	output wire auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock;
	output wire auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset;
	output wire auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock;
	output wire auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset;
	output wire auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock;
	output wire auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [1:0] monitor_io_in_a_bits_size;
	wire [7:0] monitor_io_in_a_bits_source;
	wire [20:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_size;
	wire [7:0] monitor_io_in_d_bits_source;
	wire regs_0_clock;
	wire regs_0_reset;
	wire regs_0_io_d;
	wire regs_0_io_q;
	wire regs_0_io_en;
	wire regs_1_clock;
	wire regs_1_reset;
	wire regs_1_io_d;
	wire regs_1_io_q;
	wire regs_1_io_en;
	wire regs_2_clock;
	wire regs_2_reset;
	wire regs_2_io_d;
	wire regs_2_io_q;
	wire regs_2_io_en;
	wire regs_3_clock;
	wire regs_3_reset;
	wire regs_3_io_d;
	wire regs_3_io_q;
	wire regs_3_io_en;
	wire regs_4_clock;
	wire regs_4_reset;
	wire regs_4_io_d;
	wire regs_4_io_q;
	wire regs_4_io_en;
	wire in_bits_read = auto_tile_clock_gater_in_1_a_bits_opcode == 3'h4;
	wire [9:0] in_bits_index = auto_tile_clock_gater_in_1_a_bits_address[11:2];
	wire [9:0] out_findex = in_bits_index & 10'h3f8;
	wire _out_T = out_findex == 10'h000;
	wire [7:0] _out_frontMask_T_5 = (auto_tile_clock_gater_in_1_a_bits_mask[0] ? 8'hff : 8'h00);
	wire [7:0] _out_frontMask_T_7 = (auto_tile_clock_gater_in_1_a_bits_mask[1] ? 8'hff : 8'h00);
	wire [7:0] _out_frontMask_T_9 = (auto_tile_clock_gater_in_1_a_bits_mask[2] ? 8'hff : 8'h00);
	wire [7:0] _out_frontMask_T_11 = (auto_tile_clock_gater_in_1_a_bits_mask[3] ? 8'hff : 8'h00);
	wire [31:0] out_frontMask = {_out_frontMask_T_11, _out_frontMask_T_9, _out_frontMask_T_7, _out_frontMask_T_5};
	wire out_wimask = &out_frontMask[0];
	wire [2:0] out_oindex = {in_bits_index[2], in_bits_index[1], in_bits_index[0]};
	wire [7:0] _out_frontSel_T = 8'h01 << out_oindex;
	wire out_frontSel_0 = _out_frontSel_T[0];
	wire out_wivalid_0 = (((auto_tile_clock_gater_in_1_a_valid & auto_tile_clock_gater_in_1_d_ready) & ~in_bits_read) & out_frontSel_0) & (out_findex == 10'h000);
	wire _out_T_15 = regs_0_io_q;
	wire out_frontSel_1 = _out_frontSel_T[1];
	wire out_wivalid_1 = (((auto_tile_clock_gater_in_1_a_valid & auto_tile_clock_gater_in_1_d_ready) & ~in_bits_read) & out_frontSel_1) & (out_findex == 10'h000);
	wire _out_T_22 = regs_1_io_q;
	wire out_frontSel_2 = _out_frontSel_T[2];
	wire out_wivalid_2 = (((auto_tile_clock_gater_in_1_a_valid & auto_tile_clock_gater_in_1_d_ready) & ~in_bits_read) & out_frontSel_2) & (out_findex == 10'h000);
	wire _out_T_29 = regs_2_io_q;
	wire out_frontSel_3 = _out_frontSel_T[3];
	wire out_wivalid_3 = (((auto_tile_clock_gater_in_1_a_valid & auto_tile_clock_gater_in_1_d_ready) & ~in_bits_read) & out_frontSel_3) & (out_findex == 10'h000);
	wire _out_T_36 = regs_3_io_q;
	wire out_frontSel_4 = _out_frontSel_T[4];
	wire out_wivalid_4 = (((auto_tile_clock_gater_in_1_a_valid & auto_tile_clock_gater_in_1_d_ready) & ~in_bits_read) & out_frontSel_4) & (out_findex == 10'h000);
	wire _out_T_43 = regs_4_io_q;
	wire _GEN_33 = (3'h1 == out_oindex ? _out_T : _out_T);
	wire _GEN_34 = (3'h2 == out_oindex ? _out_T : _GEN_33);
	wire _GEN_35 = (3'h3 == out_oindex ? _out_T : _GEN_34);
	wire _GEN_36 = (3'h4 == out_oindex ? _out_T : _GEN_35);
	wire _GEN_39 = (3'h7 == out_oindex) | ((3'h6 == out_oindex) | ((3'h5 == out_oindex) | _GEN_36));
	wire _GEN_41 = (3'h1 == out_oindex ? _out_T_22 : _out_T_15);
	wire _GEN_42 = (3'h2 == out_oindex ? _out_T_29 : _GEN_41);
	wire _GEN_43 = (3'h3 == out_oindex ? _out_T_36 : _GEN_42);
	wire _GEN_44 = (3'h4 == out_oindex ? _out_T_43 : _GEN_43);
	wire _GEN_45 = (3'h5 == out_oindex ? 1'h0 : _GEN_44);
	wire _GEN_46 = (3'h6 == out_oindex ? 1'h0 : _GEN_45);
	wire _GEN_47 = (3'h7 == out_oindex ? 1'h0 : _GEN_46);
	wire _out_out_bits_data_T_4 = _GEN_39 & _GEN_47;
	TLMonitor_47 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	AsyncResetRegVec_w1_i1 regs_0(
		.clock(regs_0_clock),
		.reset(regs_0_reset),
		.io_d(regs_0_io_d),
		.io_q(regs_0_io_q),
		.io_en(regs_0_io_en)
	);
	AsyncResetRegVec_w1_i1 regs_1(
		.clock(regs_1_clock),
		.reset(regs_1_reset),
		.io_d(regs_1_io_d),
		.io_q(regs_1_io_q),
		.io_en(regs_1_io_en)
	);
	AsyncResetRegVec_w1_i1 regs_2(
		.clock(regs_2_clock),
		.reset(regs_2_reset),
		.io_d(regs_2_io_d),
		.io_q(regs_2_io_q),
		.io_en(regs_2_io_en)
	);
	AsyncResetRegVec_w1_i1 regs_3(
		.clock(regs_3_clock),
		.reset(regs_3_reset),
		.io_d(regs_3_io_d),
		.io_q(regs_3_io_q),
		.io_en(regs_3_io_en)
	);
	AsyncResetRegVec_w1_i1 regs_4(
		.clock(regs_4_clock),
		.reset(regs_4_reset),
		.io_d(regs_4_io_d),
		.io_q(regs_4_io_q),
		.io_en(regs_4_io_en)
	);
	assign auto_tile_clock_gater_in_1_a_ready = auto_tile_clock_gater_in_1_d_ready;
	assign auto_tile_clock_gater_in_1_d_valid = auto_tile_clock_gater_in_1_a_valid;
	assign auto_tile_clock_gater_in_1_d_bits_opcode = {2'd0, in_bits_read};
	assign auto_tile_clock_gater_in_1_d_bits_size = auto_tile_clock_gater_in_1_a_bits_size;
	assign auto_tile_clock_gater_in_1_d_bits_source = auto_tile_clock_gater_in_1_a_bits_source;
	assign auto_tile_clock_gater_in_1_d_bits_data = {31'd0, _out_out_bits_data_T_4};
	assign auto_tile_clock_gater_out_member_allClocks_implicit_clock_clock = auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_clock;
	assign auto_tile_clock_gater_out_member_allClocks_implicit_clock_reset = auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_reset;
	assign auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock = auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_clock;
	assign auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset = auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_reset;
	assign auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock = auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_clock;
	assign auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset = auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_reset;
	assign auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock = auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_clock;
	assign auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset = auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_reset;
	assign auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock = auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_clock;
	assign auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset = auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_reset;
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_tile_clock_gater_in_1_d_ready;
	assign monitor_io_in_a_valid = auto_tile_clock_gater_in_1_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_tile_clock_gater_in_1_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_tile_clock_gater_in_1_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_tile_clock_gater_in_1_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_tile_clock_gater_in_1_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_tile_clock_gater_in_1_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_tile_clock_gater_in_1_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_tile_clock_gater_in_1_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_tile_clock_gater_in_1_d_ready;
	assign monitor_io_in_d_valid = auto_tile_clock_gater_in_1_a_valid;
	assign monitor_io_in_d_bits_opcode = {2'd0, in_bits_read};
	assign monitor_io_in_d_bits_size = auto_tile_clock_gater_in_1_a_bits_size;
	assign monitor_io_in_d_bits_source = auto_tile_clock_gater_in_1_a_bits_source;
	assign regs_0_clock = clock;
	assign regs_0_reset = auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_reset;
	assign regs_0_io_d = auto_tile_clock_gater_in_1_a_bits_data[0];
	assign regs_0_io_en = out_wivalid_0 & out_wimask;
	assign regs_1_clock = clock;
	assign regs_1_reset = auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_reset;
	assign regs_1_io_d = auto_tile_clock_gater_in_1_a_bits_data[0];
	assign regs_1_io_en = out_wivalid_1 & out_wimask;
	assign regs_2_clock = clock;
	assign regs_2_reset = auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_reset;
	assign regs_2_io_d = auto_tile_clock_gater_in_1_a_bits_data[0];
	assign regs_2_io_en = out_wivalid_2 & out_wimask;
	assign regs_3_clock = clock;
	assign regs_3_reset = auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_reset;
	assign regs_3_io_d = auto_tile_clock_gater_in_1_a_bits_data[0];
	assign regs_3_io_en = out_wivalid_3 & out_wimask;
	assign regs_4_clock = clock;
	assign regs_4_reset = auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_reset;
	assign regs_4_io_d = auto_tile_clock_gater_in_1_a_bits_data[0];
	assign regs_4_io_en = out_wivalid_4 & out_wimask;
endmodule
module TLMonitor_48 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_param,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_a_bits_corrupt,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_size,
	io_in_d_bits_source
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [2:0] io_in_a_bits_param;
	input [1:0] io_in_a_bits_size;
	input [7:0] io_in_a_bits_source;
	input [20:0] io_in_a_bits_address;
	input [3:0] io_in_a_bits_mask;
	input io_in_a_bits_corrupt;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_size;
	input [7:0] io_in_d_bits_source;
	wire [31:0] plusarg_reader_out;
	wire [31:0] plusarg_reader_1_out;
	wire _T_2 = ~reset;
	wire _source_ok_T_4 = io_in_a_bits_source <= 8'h9f;
	wire [4:0] _is_aligned_mask_T_1 = 5'h03 << io_in_a_bits_size;
	wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0];
	wire [20:0] _GEN_71 = {19'd0, is_aligned_mask};
	wire [20:0] _is_aligned_T = io_in_a_bits_address & _GEN_71;
	wire is_aligned = _is_aligned_T == 21'h000000;
	wire mask_sizeOH_shiftAmount = io_in_a_bits_size[0];
	wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount;
	wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1;
	wire _mask_T = io_in_a_bits_size >= 2'h2;
	wire mask_size = mask_sizeOH[1];
	wire mask_bit = io_in_a_bits_address[1];
	wire mask_nbit = ~mask_bit;
	wire mask_acc = _mask_T | (mask_size & mask_nbit);
	wire mask_acc_1 = _mask_T | (mask_size & mask_bit);
	wire mask_size_1 = mask_sizeOH[0];
	wire mask_bit_1 = io_in_a_bits_address[0];
	wire mask_nbit_1 = ~mask_bit_1;
	wire mask_eq_2 = mask_nbit & mask_nbit_1;
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = mask_nbit & mask_bit_1;
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = mask_bit & mask_nbit_1;
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = mask_bit & mask_bit_1;
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [3:0] mask = {mask_acc_5, mask_acc_4, mask_acc_3, mask_acc_2};
	wire _T_10 = ~_source_ok_T_4;
	wire _T_20 = io_in_a_bits_opcode == 3'h6;
	wire [20:0] _T_33 = io_in_a_bits_address ^ 21'h110000;
	wire [21:0] _T_34 = {1'b0, $signed(_T_33)};
	wire [21:0] _T_36 = $signed(_T_34) & -22'sh001000;
	wire _T_37 = $signed(_T_36) == 22'sh000000;
	wire _T_69 = io_in_a_bits_param <= 3'h2;
	wire [3:0] _T_73 = ~io_in_a_bits_mask;
	wire _T_74 = _T_73 == 4'h0;
	wire _T_78 = ~io_in_a_bits_corrupt;
	wire _T_82 = io_in_a_bits_opcode == 3'h7;
	wire _T_135 = io_in_a_bits_param != 3'h0;
	wire _T_148 = io_in_a_bits_opcode == 3'h4;
	wire _T_164 = io_in_a_bits_size <= 2'h2;
	wire _T_172 = _T_164 & _T_37;
	wire _T_183 = io_in_a_bits_param == 3'h0;
	wire _T_187 = io_in_a_bits_mask == mask;
	wire _T_195 = io_in_a_bits_opcode == 3'h0;
	wire _T_218 = _source_ok_T_4 & _T_172;
	wire _T_236 = io_in_a_bits_opcode == 3'h1;
	wire [3:0] _T_273 = ~mask;
	wire [3:0] _T_274 = io_in_a_bits_mask & _T_273;
	wire _T_275 = _T_274 == 4'h0;
	wire _T_279 = io_in_a_bits_opcode == 3'h2;
	wire _T_309 = io_in_a_bits_param <= 3'h4;
	wire _T_317 = io_in_a_bits_opcode == 3'h3;
	wire _T_347 = io_in_a_bits_param <= 3'h3;
	wire _T_355 = io_in_a_bits_opcode == 3'h5;
	wire _T_385 = io_in_a_bits_param <= 3'h1;
	wire _T_397 = io_in_d_bits_opcode <= 3'h6;
	wire _source_ok_T_10 = io_in_d_bits_source <= 8'h9f;
	wire _T_401 = io_in_d_bits_opcode == 3'h6;
	wire _T_405 = io_in_d_bits_size >= 2'h2;
	wire _T_421 = io_in_d_bits_opcode == 3'h4;
	wire _T_449 = io_in_d_bits_opcode == 3'h5;
	wire _T_478 = io_in_d_bits_opcode == 3'h0;
	wire _T_495 = io_in_d_bits_opcode == 3'h1;
	wire _T_513 = io_in_d_bits_opcode == 3'h2;
	wire a_first_done = io_in_a_ready & io_in_a_valid;
	reg a_first_counter;
	wire a_first_counter1 = a_first_counter - 1'h1;
	wire a_first = ~a_first_counter;
	reg [2:0] opcode;
	reg [2:0] param;
	reg [1:0] size;
	reg [7:0] source;
	reg [20:0] address;
	wire _T_543 = io_in_a_valid & ~a_first;
	wire _T_544 = io_in_a_bits_opcode == opcode;
	wire _T_548 = io_in_a_bits_param == param;
	wire _T_552 = io_in_a_bits_size == size;
	wire _T_556 = io_in_a_bits_source == source;
	wire _T_560 = io_in_a_bits_address == address;
	wire d_first_done = io_in_d_ready & io_in_d_valid;
	reg d_first_counter;
	wire d_first_counter1 = d_first_counter - 1'h1;
	wire d_first = ~d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] size_1;
	reg [7:0] source_1;
	wire _T_567 = io_in_d_valid & ~d_first;
	wire _T_568 = io_in_d_bits_opcode == opcode_1;
	wire _T_576 = io_in_d_bits_size == size_1;
	wire _T_580 = io_in_d_bits_source == source_1;
	reg [159:0] inflight;
	reg [639:0] inflight_opcodes;
	reg [639:0] inflight_sizes;
	reg a_first_counter_1;
	wire a_first_counter1_1 = a_first_counter_1 - 1'h1;
	wire a_first_1 = ~a_first_counter_1;
	reg d_first_counter_1;
	wire d_first_counter1_1 = d_first_counter_1 - 1'h1;
	wire d_first_1 = ~d_first_counter_1;
	wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0};
	wire [10:0] _a_opcode_lookup_T = {1'd0, _GEN_72};
	wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T;
	wire [15:0] _a_opcode_lookup_T_5 = 16'h0010 - 16'h0001;
	wire [639:0] _GEN_73 = {624'd0, _a_opcode_lookup_T_5};
	wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73;
	wire [639:0] _a_opcode_lookup_T_7 = {1'd0, _a_opcode_lookup_T_6[639:1]};
	wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T;
	wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73;
	wire [639:0] _a_size_lookup_T_7 = {1'd0, _a_size_lookup_T_6[639:1]};
	wire _T_594 = io_in_a_valid & a_first_1;
	wire [255:0] _a_set_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_a_bits_source;
	wire _T_597 = a_first_done & a_first_1;
	wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0};
	wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1;
	wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0};
	wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1;
	wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0};
	wire [10:0] _a_opcodes_set_T = {1'd0, _GEN_78};
	wire [3:0] a_opcodes_set_interm = (a_first_done & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0);
	wire [2050:0] _GEN_1 = {2047'd0, a_opcodes_set_interm};
	wire [2050:0] _a_opcodes_set_T_1 = _GEN_1 << _a_opcodes_set_T;
	wire [2:0] a_sizes_set_interm = (a_first_done & a_first_1 ? _a_sizes_set_interm_T_1 : 3'h0);
	wire [2049:0] _GEN_2 = {2047'd0, a_sizes_set_interm};
	wire [2049:0] _a_sizes_set_T_1 = _GEN_2 << _a_opcodes_set_T;
	wire [159:0] _T_599 = inflight >> io_in_a_bits_source;
	wire _T_601 = ~_T_599[0];
	wire [255:0] _GEN_16 = (a_first_done & a_first_1 ? _a_set_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2050:0] _GEN_19 = (a_first_done & a_first_1 ? _a_opcodes_set_T_1 : 2051'h0);
	wire [2049:0] _GEN_20 = (a_first_done & a_first_1 ? _a_sizes_set_T_1 : 2050'h0);
	wire _T_605 = io_in_d_valid & d_first_1;
	wire _T_607 = ~_T_401;
	wire _T_608 = (io_in_d_valid & d_first_1) & ~_T_401;
	wire [255:0] _d_clr_wo_ready_T = 256'h0000000000000000000000000000000000000000000000000000000000000001 << io_in_d_bits_source;
	wire [2062:0] _GEN_3 = {2047'd0, _a_opcode_lookup_T_5};
	wire [2062:0] _d_opcodes_clr_T_5 = _GEN_3 << _a_opcode_lookup_T;
	wire [255:0] _GEN_22 = ((d_first_done & d_first_1) & _T_607 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_23 = ((d_first_done & d_first_1) & _T_607 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source;
	wire same_cycle_resp = _T_594 & (io_in_a_bits_source == io_in_d_bits_source);
	wire [159:0] _T_618 = inflight >> io_in_d_bits_source;
	wire _T_620 = _T_618[0] | same_cycle_resp;
	wire [2:0] _GEN_27 = (3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0);
	wire [2:0] _GEN_28 = (3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27);
	wire [2:0] _GEN_29 = (3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28);
	wire [2:0] _GEN_30 = (3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29);
	wire [2:0] _GEN_31 = (3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30);
	wire [2:0] _GEN_32 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31);
	wire [2:0] _GEN_39 = (3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30);
	wire [2:0] _GEN_40 = (3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39);
	wire _T_625 = io_in_d_bits_opcode == _GEN_40;
	wire _T_626 = (io_in_d_bits_opcode == _GEN_32) | _T_625;
	wire _T_630 = io_in_a_bits_size == io_in_d_bits_size;
	wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
	wire [2:0] _GEN_43 = (3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0);
	wire [2:0] _GEN_44 = (3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43);
	wire [2:0] _GEN_45 = (3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44);
	wire [2:0] _GEN_46 = (3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45);
	wire [2:0] _GEN_47 = (3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46);
	wire [2:0] _GEN_48 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47);
	wire [2:0] _GEN_55 = (3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46);
	wire [2:0] _GEN_56 = (3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55);
	wire _T_637 = io_in_d_bits_opcode == _GEN_56;
	wire _T_638 = (io_in_d_bits_opcode == _GEN_48) | _T_637;
	wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
	wire [3:0] _GEN_82 = {2'd0, io_in_d_bits_size};
	wire _T_642 = _GEN_82 == a_size_lookup;
	wire _T_652 = (((_T_605 & a_first_1) & io_in_a_valid) & _same_cycle_resp_T_2) & _T_607;
	wire _T_654 = ~io_in_d_ready | io_in_a_ready;
	wire [159:0] a_set = _GEN_16[159:0];
	wire [159:0] _inflight_T = inflight | a_set;
	wire [159:0] d_clr = _GEN_22[159:0];
	wire [159:0] _inflight_T_1 = ~d_clr;
	wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1;
	wire [639:0] a_opcodes_set = _GEN_19[639:0];
	wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set;
	wire [639:0] d_opcodes_clr = _GEN_23[639:0];
	wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr;
	wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1;
	wire [639:0] a_sizes_set = _GEN_20[639:0];
	wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set;
	wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1;
	reg [31:0] watchdog;
	wire _T_663 = (~(|inflight) | (plusarg_reader_out == 32'h00000000)) | (watchdog < plusarg_reader_out);
	wire [31:0] _watchdog_T_1 = watchdog + 32'h00000001;
	reg [159:0] inflight_1;
	reg [639:0] inflight_sizes_1;
	reg d_first_counter_2;
	wire d_first_counter1_2 = d_first_counter_2 - 1'h1;
	wire d_first_2 = ~d_first_counter_2;
	wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T;
	wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73;
	wire [639:0] _c_size_lookup_T_7 = {1'd0, _c_size_lookup_T_6[639:1]};
	wire _T_689 = (io_in_d_valid & d_first_2) & _T_401;
	wire [255:0] _GEN_67 = ((d_first_done & d_first_2) & _T_401 ? _d_clr_wo_ready_T : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	wire [2062:0] _GEN_68 = ((d_first_done & d_first_2) & _T_401 ? _d_opcodes_clr_T_5 : 2063'h0);
	wire [159:0] _T_697 = inflight_1 >> io_in_d_bits_source;
	wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
	wire _T_707 = _GEN_82 == c_size_lookup;
	wire [159:0] d_clr_1 = _GEN_67[159:0];
	wire [159:0] _inflight_T_4 = ~d_clr_1;
	wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4;
	wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0];
	wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1;
	wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4;
	reg [31:0] watchdog_1;
	wire _T_727 = (~(|inflight_1) | (plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < plusarg_reader_1_out);
	wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h00000001;
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader(.out(plusarg_reader_out));
	plusarg_reader #(
		.FORMAT("tilelink_timeout=%d"),
		.DEFAULT(0),
		.WIDTH(32)
	) plusarg_reader_1(.out(plusarg_reader_1_out));
	always @(posedge clock) begin
		if (reset)
			a_first_counter <= 1'h0;
		else if (a_first_done)
			if (a_first)
				a_first_counter <= 1'h0;
			else
				a_first_counter <= a_first_counter1;
		if (a_first_done & a_first)
			opcode <= io_in_a_bits_opcode;
		if (a_first_done & a_first)
			param <= io_in_a_bits_param;
		if (a_first_done & a_first)
			size <= io_in_a_bits_size;
		if (a_first_done & a_first)
			source <= io_in_a_bits_source;
		if (a_first_done & a_first)
			address <= io_in_a_bits_address;
		if (reset)
			d_first_counter <= 1'h0;
		else if (d_first_done)
			if (d_first)
				d_first_counter <= 1'h0;
			else
				d_first_counter <= d_first_counter1;
		if (d_first_done & d_first)
			opcode_1 <= io_in_d_bits_opcode;
		if (d_first_done & d_first)
			size_1 <= io_in_d_bits_size;
		if (d_first_done & d_first)
			source_1 <= io_in_d_bits_source;
		if (reset)
			inflight <= 160'h0000000000000000000000000000000000000000;
		else
			inflight <= _inflight_T_2;
		if (reset)
			inflight_opcodes <= 640'h0;
		else
			inflight_opcodes <= _inflight_opcodes_T_2;
		if (reset)
			inflight_sizes <= 640'h0;
		else
			inflight_sizes <= _inflight_sizes_T_2;
		if (reset)
			a_first_counter_1 <= 1'h0;
		else if (a_first_done)
			if (a_first_1)
				a_first_counter_1 <= 1'h0;
			else
				a_first_counter_1 <= a_first_counter1_1;
		if (reset)
			d_first_counter_1 <= 1'h0;
		else if (d_first_done)
			if (d_first_1)
				d_first_counter_1 <= 1'h0;
			else
				d_first_counter_1 <= d_first_counter1_1;
		if (reset)
			watchdog <= 32'h00000000;
		else if (a_first_done | d_first_done)
			watchdog <= 32'h00000000;
		else
			watchdog <= _watchdog_T_1;
		if (reset)
			inflight_1 <= 160'h0000000000000000000000000000000000000000;
		else
			inflight_1 <= _inflight_T_5;
		if (reset)
			inflight_sizes_1 <= 640'h0;
		else
			inflight_sizes_1 <= _inflight_sizes_T_5;
		if (reset)
			d_first_counter_2 <= 1'h0;
		else if (d_first_done)
			if (d_first_2)
				d_first_counter_2 <= 1'h0;
			else
				d_first_counter_2 <= d_first_counter1_2;
		if (reset)
			watchdog_1 <= 32'h00000000;
		else if (d_first_done)
			watchdog_1 <= 32'h00000000;
		else
			watchdog_1 <= _watchdog_T_3;
	end
endmodule
module AsyncResetRegVec_w1_i0_5 (
	clock,
	reset,
	io_d,
	io_q,
	io_en
);
	input clock;
	input reset;
	input io_d;
	output wire io_q;
	input io_en;
	reg reg_;
	assign io_q = reg_;
	always @(posedge clock or posedge reset)
		if (reset)
			reg_ <= 1'h0;
		else if (io_en)
			reg_ <= io_d;
endmodule
module TileResetSetter (
	clock,
	reset,
	auto_clock_in_member_allClocks_implicit_clock_clock,
	auto_clock_in_member_allClocks_implicit_clock_reset,
	auto_clock_in_member_allClocks_subsystem_cbus_0_clock,
	auto_clock_in_member_allClocks_subsystem_cbus_0_reset,
	auto_clock_in_member_allClocks_subsystem_fbus_0_clock,
	auto_clock_in_member_allClocks_subsystem_fbus_0_reset,
	auto_clock_in_member_allClocks_subsystem_pbus_0_clock,
	auto_clock_in_member_allClocks_subsystem_pbus_0_reset,
	auto_clock_in_member_allClocks_subsystem_sbus_0_clock,
	auto_clock_in_member_allClocks_subsystem_sbus_0_reset,
	auto_clock_out_member_allClocks_implicit_clock_clock,
	auto_clock_out_member_allClocks_implicit_clock_reset,
	auto_clock_out_member_allClocks_subsystem_cbus_0_clock,
	auto_clock_out_member_allClocks_subsystem_cbus_0_reset,
	auto_clock_out_member_allClocks_subsystem_fbus_0_clock,
	auto_clock_out_member_allClocks_subsystem_fbus_0_reset,
	auto_clock_out_member_allClocks_subsystem_pbus_0_clock,
	auto_clock_out_member_allClocks_subsystem_pbus_0_reset,
	auto_clock_out_member_allClocks_subsystem_sbus_0_clock,
	auto_clock_out_member_allClocks_subsystem_sbus_0_reset,
	auto_tl_in_a_ready,
	auto_tl_in_a_valid,
	auto_tl_in_a_bits_opcode,
	auto_tl_in_a_bits_param,
	auto_tl_in_a_bits_size,
	auto_tl_in_a_bits_source,
	auto_tl_in_a_bits_address,
	auto_tl_in_a_bits_mask,
	auto_tl_in_a_bits_data,
	auto_tl_in_a_bits_corrupt,
	auto_tl_in_d_ready,
	auto_tl_in_d_valid,
	auto_tl_in_d_bits_opcode,
	auto_tl_in_d_bits_size,
	auto_tl_in_d_bits_source,
	auto_tl_in_d_bits_data
);
	input clock;
	input reset;
	input auto_clock_in_member_allClocks_implicit_clock_clock;
	input auto_clock_in_member_allClocks_implicit_clock_reset;
	input auto_clock_in_member_allClocks_subsystem_cbus_0_clock;
	input auto_clock_in_member_allClocks_subsystem_cbus_0_reset;
	input auto_clock_in_member_allClocks_subsystem_fbus_0_clock;
	input auto_clock_in_member_allClocks_subsystem_fbus_0_reset;
	input auto_clock_in_member_allClocks_subsystem_pbus_0_clock;
	input auto_clock_in_member_allClocks_subsystem_pbus_0_reset;
	input auto_clock_in_member_allClocks_subsystem_sbus_0_clock;
	input auto_clock_in_member_allClocks_subsystem_sbus_0_reset;
	output wire auto_clock_out_member_allClocks_implicit_clock_clock;
	output wire auto_clock_out_member_allClocks_implicit_clock_reset;
	output wire auto_clock_out_member_allClocks_subsystem_cbus_0_clock;
	output wire auto_clock_out_member_allClocks_subsystem_cbus_0_reset;
	output wire auto_clock_out_member_allClocks_subsystem_fbus_0_clock;
	output wire auto_clock_out_member_allClocks_subsystem_fbus_0_reset;
	output wire auto_clock_out_member_allClocks_subsystem_pbus_0_clock;
	output wire auto_clock_out_member_allClocks_subsystem_pbus_0_reset;
	output wire auto_clock_out_member_allClocks_subsystem_sbus_0_clock;
	output wire auto_clock_out_member_allClocks_subsystem_sbus_0_reset;
	output wire auto_tl_in_a_ready;
	input auto_tl_in_a_valid;
	input [2:0] auto_tl_in_a_bits_opcode;
	input [2:0] auto_tl_in_a_bits_param;
	input [1:0] auto_tl_in_a_bits_size;
	input [7:0] auto_tl_in_a_bits_source;
	input [20:0] auto_tl_in_a_bits_address;
	input [3:0] auto_tl_in_a_bits_mask;
	input [31:0] auto_tl_in_a_bits_data;
	input auto_tl_in_a_bits_corrupt;
	input auto_tl_in_d_ready;
	output wire auto_tl_in_d_valid;
	output wire [2:0] auto_tl_in_d_bits_opcode;
	output wire [1:0] auto_tl_in_d_bits_size;
	output wire [7:0] auto_tl_in_d_bits_source;
	output wire [31:0] auto_tl_in_d_bits_data;
	wire monitor_clock;
	wire monitor_reset;
	wire monitor_io_in_a_ready;
	wire monitor_io_in_a_valid;
	wire [2:0] monitor_io_in_a_bits_opcode;
	wire [2:0] monitor_io_in_a_bits_param;
	wire [1:0] monitor_io_in_a_bits_size;
	wire [7:0] monitor_io_in_a_bits_source;
	wire [20:0] monitor_io_in_a_bits_address;
	wire [3:0] monitor_io_in_a_bits_mask;
	wire monitor_io_in_a_bits_corrupt;
	wire monitor_io_in_d_ready;
	wire monitor_io_in_d_valid;
	wire [2:0] monitor_io_in_d_bits_opcode;
	wire [1:0] monitor_io_in_d_bits_size;
	wire [7:0] monitor_io_in_d_bits_source;
	wire r_tile_resets_0_clock;
	wire r_tile_resets_0_reset;
	wire r_tile_resets_0_io_d;
	wire r_tile_resets_0_io_q;
	wire r_tile_resets_0_io_en;
	wire in_bits_read = auto_tl_in_a_bits_opcode == 3'h4;
	wire [9:0] in_bits_index = auto_tl_in_a_bits_address[11:2];
	wire [7:0] _out_frontMask_T_5 = (auto_tl_in_a_bits_mask[0] ? 8'hff : 8'h00);
	wire [7:0] _out_frontMask_T_7 = (auto_tl_in_a_bits_mask[1] ? 8'hff : 8'h00);
	wire [7:0] _out_frontMask_T_9 = (auto_tl_in_a_bits_mask[2] ? 8'hff : 8'h00);
	wire [7:0] _out_frontMask_T_11 = (auto_tl_in_a_bits_mask[3] ? 8'hff : 8'h00);
	wire [31:0] out_frontMask = {_out_frontMask_T_11, _out_frontMask_T_9, _out_frontMask_T_7, _out_frontMask_T_5};
	wire out_wimask = &out_frontMask[0];
	wire out_wivalid_0 = ((auto_tl_in_a_valid & auto_tl_in_d_ready) & ~in_bits_read) & (in_bits_index == 10'h000);
	wire _out_out_bits_data_T_4 = (in_bits_index == 10'h000) & r_tile_resets_0_io_q;
	TLMonitor_48 monitor(
		.clock(monitor_clock),
		.reset(monitor_reset),
		.io_in_a_ready(monitor_io_in_a_ready),
		.io_in_a_valid(monitor_io_in_a_valid),
		.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
		.io_in_a_bits_param(monitor_io_in_a_bits_param),
		.io_in_a_bits_size(monitor_io_in_a_bits_size),
		.io_in_a_bits_source(monitor_io_in_a_bits_source),
		.io_in_a_bits_address(monitor_io_in_a_bits_address),
		.io_in_a_bits_mask(monitor_io_in_a_bits_mask),
		.io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
		.io_in_d_ready(monitor_io_in_d_ready),
		.io_in_d_valid(monitor_io_in_d_valid),
		.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
		.io_in_d_bits_size(monitor_io_in_d_bits_size),
		.io_in_d_bits_source(monitor_io_in_d_bits_source)
	);
	AsyncResetRegVec_w1_i0_5 r_tile_resets_0(
		.clock(r_tile_resets_0_clock),
		.reset(r_tile_resets_0_reset),
		.io_d(r_tile_resets_0_io_d),
		.io_q(r_tile_resets_0_io_q),
		.io_en(r_tile_resets_0_io_en)
	);
	assign auto_clock_out_member_allClocks_implicit_clock_clock = auto_clock_in_member_allClocks_implicit_clock_clock;
	assign auto_clock_out_member_allClocks_implicit_clock_reset = auto_clock_in_member_allClocks_implicit_clock_reset;
	assign auto_clock_out_member_allClocks_subsystem_cbus_0_clock = auto_clock_in_member_allClocks_subsystem_cbus_0_clock;
	assign auto_clock_out_member_allClocks_subsystem_cbus_0_reset = auto_clock_in_member_allClocks_subsystem_cbus_0_reset;
	assign auto_clock_out_member_allClocks_subsystem_fbus_0_clock = auto_clock_in_member_allClocks_subsystem_fbus_0_clock;
	assign auto_clock_out_member_allClocks_subsystem_fbus_0_reset = auto_clock_in_member_allClocks_subsystem_fbus_0_reset;
	assign auto_clock_out_member_allClocks_subsystem_pbus_0_clock = auto_clock_in_member_allClocks_subsystem_pbus_0_clock;
	assign auto_clock_out_member_allClocks_subsystem_pbus_0_reset = auto_clock_in_member_allClocks_subsystem_pbus_0_reset;
	assign auto_clock_out_member_allClocks_subsystem_sbus_0_clock = auto_clock_in_member_allClocks_subsystem_sbus_0_clock;
	assign auto_clock_out_member_allClocks_subsystem_sbus_0_reset = auto_clock_in_member_allClocks_subsystem_sbus_0_reset;
	assign auto_tl_in_a_ready = auto_tl_in_d_ready;
	assign auto_tl_in_d_valid = auto_tl_in_a_valid;
	assign auto_tl_in_d_bits_opcode = {2'd0, in_bits_read};
	assign auto_tl_in_d_bits_size = auto_tl_in_a_bits_size;
	assign auto_tl_in_d_bits_source = auto_tl_in_a_bits_source;
	assign auto_tl_in_d_bits_data = {31'd0, _out_out_bits_data_T_4};
	assign monitor_clock = clock;
	assign monitor_reset = reset;
	assign monitor_io_in_a_ready = auto_tl_in_d_ready;
	assign monitor_io_in_a_valid = auto_tl_in_a_valid;
	assign monitor_io_in_a_bits_opcode = auto_tl_in_a_bits_opcode;
	assign monitor_io_in_a_bits_param = auto_tl_in_a_bits_param;
	assign monitor_io_in_a_bits_size = auto_tl_in_a_bits_size;
	assign monitor_io_in_a_bits_source = auto_tl_in_a_bits_source;
	assign monitor_io_in_a_bits_address = auto_tl_in_a_bits_address;
	assign monitor_io_in_a_bits_mask = auto_tl_in_a_bits_mask;
	assign monitor_io_in_a_bits_corrupt = auto_tl_in_a_bits_corrupt;
	assign monitor_io_in_d_ready = auto_tl_in_d_ready;
	assign monitor_io_in_d_valid = auto_tl_in_a_valid;
	assign monitor_io_in_d_bits_opcode = {2'd0, in_bits_read};
	assign monitor_io_in_d_bits_size = auto_tl_in_a_bits_size;
	assign monitor_io_in_d_bits_source = auto_tl_in_a_bits_source;
	assign r_tile_resets_0_clock = clock;
	assign r_tile_resets_0_reset = 1'h1;
	assign r_tile_resets_0_io_d = auto_tl_in_a_bits_data[0];
	assign r_tile_resets_0_io_en = out_wivalid_0 & out_wimask;
endmodule
module ClockSinkDomain_4 (
	auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock,
	auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset,
	auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock,
	auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset,
	auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock,
	auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset,
	auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock,
	auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset,
	auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock,
	auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset,
	auto_tileResetSetter_tl_in_a_ready,
	auto_tileResetSetter_tl_in_a_valid,
	auto_tileResetSetter_tl_in_a_bits_opcode,
	auto_tileResetSetter_tl_in_a_bits_param,
	auto_tileResetSetter_tl_in_a_bits_size,
	auto_tileResetSetter_tl_in_a_bits_source,
	auto_tileResetSetter_tl_in_a_bits_address,
	auto_tileResetSetter_tl_in_a_bits_mask,
	auto_tileResetSetter_tl_in_a_bits_data,
	auto_tileResetSetter_tl_in_a_bits_corrupt,
	auto_tileResetSetter_tl_in_d_ready,
	auto_tileResetSetter_tl_in_d_valid,
	auto_tileResetSetter_tl_in_d_bits_opcode,
	auto_tileResetSetter_tl_in_d_bits_size,
	auto_tileResetSetter_tl_in_d_bits_source,
	auto_tileResetSetter_tl_in_d_bits_data,
	auto_tileClockGater_tile_clock_gater_in_a_ready,
	auto_tileClockGater_tile_clock_gater_in_a_valid,
	auto_tileClockGater_tile_clock_gater_in_a_bits_opcode,
	auto_tileClockGater_tile_clock_gater_in_a_bits_param,
	auto_tileClockGater_tile_clock_gater_in_a_bits_size,
	auto_tileClockGater_tile_clock_gater_in_a_bits_source,
	auto_tileClockGater_tile_clock_gater_in_a_bits_address,
	auto_tileClockGater_tile_clock_gater_in_a_bits_mask,
	auto_tileClockGater_tile_clock_gater_in_a_bits_data,
	auto_tileClockGater_tile_clock_gater_in_a_bits_corrupt,
	auto_tileClockGater_tile_clock_gater_in_d_ready,
	auto_tileClockGater_tile_clock_gater_in_d_valid,
	auto_tileClockGater_tile_clock_gater_in_d_bits_opcode,
	auto_tileClockGater_tile_clock_gater_in_d_bits_size,
	auto_tileClockGater_tile_clock_gater_in_d_bits_source,
	auto_tileClockGater_tile_clock_gater_in_d_bits_data,
	auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_clock,
	auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_reset,
	auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock,
	auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset,
	auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock,
	auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset,
	auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock,
	auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset,
	auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock,
	auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset,
	auto_clock_in_clock,
	auto_clock_in_reset
);
	input auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock;
	input auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset;
	input auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock;
	input auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset;
	input auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock;
	input auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset;
	input auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock;
	input auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset;
	input auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock;
	input auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset;
	output wire auto_tileResetSetter_tl_in_a_ready;
	input auto_tileResetSetter_tl_in_a_valid;
	input [2:0] auto_tileResetSetter_tl_in_a_bits_opcode;
	input [2:0] auto_tileResetSetter_tl_in_a_bits_param;
	input [1:0] auto_tileResetSetter_tl_in_a_bits_size;
	input [7:0] auto_tileResetSetter_tl_in_a_bits_source;
	input [20:0] auto_tileResetSetter_tl_in_a_bits_address;
	input [3:0] auto_tileResetSetter_tl_in_a_bits_mask;
	input [31:0] auto_tileResetSetter_tl_in_a_bits_data;
	input auto_tileResetSetter_tl_in_a_bits_corrupt;
	input auto_tileResetSetter_tl_in_d_ready;
	output wire auto_tileResetSetter_tl_in_d_valid;
	output wire [2:0] auto_tileResetSetter_tl_in_d_bits_opcode;
	output wire [1:0] auto_tileResetSetter_tl_in_d_bits_size;
	output wire [7:0] auto_tileResetSetter_tl_in_d_bits_source;
	output wire [31:0] auto_tileResetSetter_tl_in_d_bits_data;
	output wire auto_tileClockGater_tile_clock_gater_in_a_ready;
	input auto_tileClockGater_tile_clock_gater_in_a_valid;
	input [2:0] auto_tileClockGater_tile_clock_gater_in_a_bits_opcode;
	input [2:0] auto_tileClockGater_tile_clock_gater_in_a_bits_param;
	input [1:0] auto_tileClockGater_tile_clock_gater_in_a_bits_size;
	input [7:0] auto_tileClockGater_tile_clock_gater_in_a_bits_source;
	input [20:0] auto_tileClockGater_tile_clock_gater_in_a_bits_address;
	input [3:0] auto_tileClockGater_tile_clock_gater_in_a_bits_mask;
	input [31:0] auto_tileClockGater_tile_clock_gater_in_a_bits_data;
	input auto_tileClockGater_tile_clock_gater_in_a_bits_corrupt;
	input auto_tileClockGater_tile_clock_gater_in_d_ready;
	output wire auto_tileClockGater_tile_clock_gater_in_d_valid;
	output wire [2:0] auto_tileClockGater_tile_clock_gater_in_d_bits_opcode;
	output wire [1:0] auto_tileClockGater_tile_clock_gater_in_d_bits_size;
	output wire [7:0] auto_tileClockGater_tile_clock_gater_in_d_bits_source;
	output wire [31:0] auto_tileClockGater_tile_clock_gater_in_d_bits_data;
	output wire auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_clock;
	output wire auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_reset;
	output wire auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock;
	output wire auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset;
	output wire auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock;
	output wire auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset;
	output wire auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock;
	output wire auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset;
	output wire auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock;
	output wire auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset;
	input auto_clock_in_clock;
	input auto_clock_in_reset;
	wire tileClockGater_clock;
	wire tileClockGater_reset;
	wire tileClockGater_auto_tile_clock_gater_in_1_a_ready;
	wire tileClockGater_auto_tile_clock_gater_in_1_a_valid;
	wire [2:0] tileClockGater_auto_tile_clock_gater_in_1_a_bits_opcode;
	wire [2:0] tileClockGater_auto_tile_clock_gater_in_1_a_bits_param;
	wire [1:0] tileClockGater_auto_tile_clock_gater_in_1_a_bits_size;
	wire [7:0] tileClockGater_auto_tile_clock_gater_in_1_a_bits_source;
	wire [20:0] tileClockGater_auto_tile_clock_gater_in_1_a_bits_address;
	wire [3:0] tileClockGater_auto_tile_clock_gater_in_1_a_bits_mask;
	wire [31:0] tileClockGater_auto_tile_clock_gater_in_1_a_bits_data;
	wire tileClockGater_auto_tile_clock_gater_in_1_a_bits_corrupt;
	wire tileClockGater_auto_tile_clock_gater_in_1_d_ready;
	wire tileClockGater_auto_tile_clock_gater_in_1_d_valid;
	wire [2:0] tileClockGater_auto_tile_clock_gater_in_1_d_bits_opcode;
	wire [1:0] tileClockGater_auto_tile_clock_gater_in_1_d_bits_size;
	wire [7:0] tileClockGater_auto_tile_clock_gater_in_1_d_bits_source;
	wire [31:0] tileClockGater_auto_tile_clock_gater_in_1_d_bits_data;
	wire tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_clock;
	wire tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_reset;
	wire tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_clock;
	wire tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_reset;
	wire tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_clock;
	wire tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_reset;
	wire tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_clock;
	wire tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_reset;
	wire tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_clock;
	wire tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_reset;
	wire tileClockGater_auto_tile_clock_gater_out_member_allClocks_implicit_clock_clock;
	wire tileClockGater_auto_tile_clock_gater_out_member_allClocks_implicit_clock_reset;
	wire tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock;
	wire tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset;
	wire tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock;
	wire tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset;
	wire tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock;
	wire tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset;
	wire tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock;
	wire tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset;
	wire tileResetSetter_clock;
	wire tileResetSetter_reset;
	wire tileResetSetter_auto_clock_in_member_allClocks_implicit_clock_clock;
	wire tileResetSetter_auto_clock_in_member_allClocks_implicit_clock_reset;
	wire tileResetSetter_auto_clock_in_member_allClocks_subsystem_cbus_0_clock;
	wire tileResetSetter_auto_clock_in_member_allClocks_subsystem_cbus_0_reset;
	wire tileResetSetter_auto_clock_in_member_allClocks_subsystem_fbus_0_clock;
	wire tileResetSetter_auto_clock_in_member_allClocks_subsystem_fbus_0_reset;
	wire tileResetSetter_auto_clock_in_member_allClocks_subsystem_pbus_0_clock;
	wire tileResetSetter_auto_clock_in_member_allClocks_subsystem_pbus_0_reset;
	wire tileResetSetter_auto_clock_in_member_allClocks_subsystem_sbus_0_clock;
	wire tileResetSetter_auto_clock_in_member_allClocks_subsystem_sbus_0_reset;
	wire tileResetSetter_auto_clock_out_member_allClocks_implicit_clock_clock;
	wire tileResetSetter_auto_clock_out_member_allClocks_implicit_clock_reset;
	wire tileResetSetter_auto_clock_out_member_allClocks_subsystem_cbus_0_clock;
	wire tileResetSetter_auto_clock_out_member_allClocks_subsystem_cbus_0_reset;
	wire tileResetSetter_auto_clock_out_member_allClocks_subsystem_fbus_0_clock;
	wire tileResetSetter_auto_clock_out_member_allClocks_subsystem_fbus_0_reset;
	wire tileResetSetter_auto_clock_out_member_allClocks_subsystem_pbus_0_clock;
	wire tileResetSetter_auto_clock_out_member_allClocks_subsystem_pbus_0_reset;
	wire tileResetSetter_auto_clock_out_member_allClocks_subsystem_sbus_0_clock;
	wire tileResetSetter_auto_clock_out_member_allClocks_subsystem_sbus_0_reset;
	wire tileResetSetter_auto_tl_in_a_ready;
	wire tileResetSetter_auto_tl_in_a_valid;
	wire [2:0] tileResetSetter_auto_tl_in_a_bits_opcode;
	wire [2:0] tileResetSetter_auto_tl_in_a_bits_param;
	wire [1:0] tileResetSetter_auto_tl_in_a_bits_size;
	wire [7:0] tileResetSetter_auto_tl_in_a_bits_source;
	wire [20:0] tileResetSetter_auto_tl_in_a_bits_address;
	wire [3:0] tileResetSetter_auto_tl_in_a_bits_mask;
	wire [31:0] tileResetSetter_auto_tl_in_a_bits_data;
	wire tileResetSetter_auto_tl_in_a_bits_corrupt;
	wire tileResetSetter_auto_tl_in_d_ready;
	wire tileResetSetter_auto_tl_in_d_valid;
	wire [2:0] tileResetSetter_auto_tl_in_d_bits_opcode;
	wire [1:0] tileResetSetter_auto_tl_in_d_bits_size;
	wire [7:0] tileResetSetter_auto_tl_in_d_bits_source;
	wire [31:0] tileResetSetter_auto_tl_in_d_bits_data;
	TileClockGater tileClockGater(
		.clock(tileClockGater_clock),
		.reset(tileClockGater_reset),
		.auto_tile_clock_gater_in_1_a_ready(tileClockGater_auto_tile_clock_gater_in_1_a_ready),
		.auto_tile_clock_gater_in_1_a_valid(tileClockGater_auto_tile_clock_gater_in_1_a_valid),
		.auto_tile_clock_gater_in_1_a_bits_opcode(tileClockGater_auto_tile_clock_gater_in_1_a_bits_opcode),
		.auto_tile_clock_gater_in_1_a_bits_param(tileClockGater_auto_tile_clock_gater_in_1_a_bits_param),
		.auto_tile_clock_gater_in_1_a_bits_size(tileClockGater_auto_tile_clock_gater_in_1_a_bits_size),
		.auto_tile_clock_gater_in_1_a_bits_source(tileClockGater_auto_tile_clock_gater_in_1_a_bits_source),
		.auto_tile_clock_gater_in_1_a_bits_address(tileClockGater_auto_tile_clock_gater_in_1_a_bits_address),
		.auto_tile_clock_gater_in_1_a_bits_mask(tileClockGater_auto_tile_clock_gater_in_1_a_bits_mask),
		.auto_tile_clock_gater_in_1_a_bits_data(tileClockGater_auto_tile_clock_gater_in_1_a_bits_data),
		.auto_tile_clock_gater_in_1_a_bits_corrupt(tileClockGater_auto_tile_clock_gater_in_1_a_bits_corrupt),
		.auto_tile_clock_gater_in_1_d_ready(tileClockGater_auto_tile_clock_gater_in_1_d_ready),
		.auto_tile_clock_gater_in_1_d_valid(tileClockGater_auto_tile_clock_gater_in_1_d_valid),
		.auto_tile_clock_gater_in_1_d_bits_opcode(tileClockGater_auto_tile_clock_gater_in_1_d_bits_opcode),
		.auto_tile_clock_gater_in_1_d_bits_size(tileClockGater_auto_tile_clock_gater_in_1_d_bits_size),
		.auto_tile_clock_gater_in_1_d_bits_source(tileClockGater_auto_tile_clock_gater_in_1_d_bits_source),
		.auto_tile_clock_gater_in_1_d_bits_data(tileClockGater_auto_tile_clock_gater_in_1_d_bits_data),
		.auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_clock(tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_clock),
		.auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_reset(tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_reset),
		.auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_clock(tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_clock),
		.auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_reset(tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_reset),
		.auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_clock(tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_clock),
		.auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_reset(tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_reset),
		.auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_clock(tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_clock),
		.auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_reset(tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_reset),
		.auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_clock(tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_clock),
		.auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_reset(tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_reset),
		.auto_tile_clock_gater_out_member_allClocks_implicit_clock_clock(tileClockGater_auto_tile_clock_gater_out_member_allClocks_implicit_clock_clock),
		.auto_tile_clock_gater_out_member_allClocks_implicit_clock_reset(tileClockGater_auto_tile_clock_gater_out_member_allClocks_implicit_clock_reset),
		.auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock(tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock),
		.auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset(tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset),
		.auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock(tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock),
		.auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset(tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset),
		.auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock(tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock),
		.auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset(tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset),
		.auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock(tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock),
		.auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset(tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset)
	);
	TileResetSetter tileResetSetter(
		.clock(tileResetSetter_clock),
		.reset(tileResetSetter_reset),
		.auto_clock_in_member_allClocks_implicit_clock_clock(tileResetSetter_auto_clock_in_member_allClocks_implicit_clock_clock),
		.auto_clock_in_member_allClocks_implicit_clock_reset(tileResetSetter_auto_clock_in_member_allClocks_implicit_clock_reset),
		.auto_clock_in_member_allClocks_subsystem_cbus_0_clock(tileResetSetter_auto_clock_in_member_allClocks_subsystem_cbus_0_clock),
		.auto_clock_in_member_allClocks_subsystem_cbus_0_reset(tileResetSetter_auto_clock_in_member_allClocks_subsystem_cbus_0_reset),
		.auto_clock_in_member_allClocks_subsystem_fbus_0_clock(tileResetSetter_auto_clock_in_member_allClocks_subsystem_fbus_0_clock),
		.auto_clock_in_member_allClocks_subsystem_fbus_0_reset(tileResetSetter_auto_clock_in_member_allClocks_subsystem_fbus_0_reset),
		.auto_clock_in_member_allClocks_subsystem_pbus_0_clock(tileResetSetter_auto_clock_in_member_allClocks_subsystem_pbus_0_clock),
		.auto_clock_in_member_allClocks_subsystem_pbus_0_reset(tileResetSetter_auto_clock_in_member_allClocks_subsystem_pbus_0_reset),
		.auto_clock_in_member_allClocks_subsystem_sbus_0_clock(tileResetSetter_auto_clock_in_member_allClocks_subsystem_sbus_0_clock),
		.auto_clock_in_member_allClocks_subsystem_sbus_0_reset(tileResetSetter_auto_clock_in_member_allClocks_subsystem_sbus_0_reset),
		.auto_clock_out_member_allClocks_implicit_clock_clock(tileResetSetter_auto_clock_out_member_allClocks_implicit_clock_clock),
		.auto_clock_out_member_allClocks_implicit_clock_reset(tileResetSetter_auto_clock_out_member_allClocks_implicit_clock_reset),
		.auto_clock_out_member_allClocks_subsystem_cbus_0_clock(tileResetSetter_auto_clock_out_member_allClocks_subsystem_cbus_0_clock),
		.auto_clock_out_member_allClocks_subsystem_cbus_0_reset(tileResetSetter_auto_clock_out_member_allClocks_subsystem_cbus_0_reset),
		.auto_clock_out_member_allClocks_subsystem_fbus_0_clock(tileResetSetter_auto_clock_out_member_allClocks_subsystem_fbus_0_clock),
		.auto_clock_out_member_allClocks_subsystem_fbus_0_reset(tileResetSetter_auto_clock_out_member_allClocks_subsystem_fbus_0_reset),
		.auto_clock_out_member_allClocks_subsystem_pbus_0_clock(tileResetSetter_auto_clock_out_member_allClocks_subsystem_pbus_0_clock),
		.auto_clock_out_member_allClocks_subsystem_pbus_0_reset(tileResetSetter_auto_clock_out_member_allClocks_subsystem_pbus_0_reset),
		.auto_clock_out_member_allClocks_subsystem_sbus_0_clock(tileResetSetter_auto_clock_out_member_allClocks_subsystem_sbus_0_clock),
		.auto_clock_out_member_allClocks_subsystem_sbus_0_reset(tileResetSetter_auto_clock_out_member_allClocks_subsystem_sbus_0_reset),
		.auto_tl_in_a_ready(tileResetSetter_auto_tl_in_a_ready),
		.auto_tl_in_a_valid(tileResetSetter_auto_tl_in_a_valid),
		.auto_tl_in_a_bits_opcode(tileResetSetter_auto_tl_in_a_bits_opcode),
		.auto_tl_in_a_bits_param(tileResetSetter_auto_tl_in_a_bits_param),
		.auto_tl_in_a_bits_size(tileResetSetter_auto_tl_in_a_bits_size),
		.auto_tl_in_a_bits_source(tileResetSetter_auto_tl_in_a_bits_source),
		.auto_tl_in_a_bits_address(tileResetSetter_auto_tl_in_a_bits_address),
		.auto_tl_in_a_bits_mask(tileResetSetter_auto_tl_in_a_bits_mask),
		.auto_tl_in_a_bits_data(tileResetSetter_auto_tl_in_a_bits_data),
		.auto_tl_in_a_bits_corrupt(tileResetSetter_auto_tl_in_a_bits_corrupt),
		.auto_tl_in_d_ready(tileResetSetter_auto_tl_in_d_ready),
		.auto_tl_in_d_valid(tileResetSetter_auto_tl_in_d_valid),
		.auto_tl_in_d_bits_opcode(tileResetSetter_auto_tl_in_d_bits_opcode),
		.auto_tl_in_d_bits_size(tileResetSetter_auto_tl_in_d_bits_size),
		.auto_tl_in_d_bits_source(tileResetSetter_auto_tl_in_d_bits_source),
		.auto_tl_in_d_bits_data(tileResetSetter_auto_tl_in_d_bits_data)
	);
	assign auto_tileResetSetter_tl_in_a_ready = tileResetSetter_auto_tl_in_a_ready;
	assign auto_tileResetSetter_tl_in_d_valid = tileResetSetter_auto_tl_in_d_valid;
	assign auto_tileResetSetter_tl_in_d_bits_opcode = tileResetSetter_auto_tl_in_d_bits_opcode;
	assign auto_tileResetSetter_tl_in_d_bits_size = tileResetSetter_auto_tl_in_d_bits_size;
	assign auto_tileResetSetter_tl_in_d_bits_source = tileResetSetter_auto_tl_in_d_bits_source;
	assign auto_tileResetSetter_tl_in_d_bits_data = tileResetSetter_auto_tl_in_d_bits_data;
	assign auto_tileClockGater_tile_clock_gater_in_a_ready = tileClockGater_auto_tile_clock_gater_in_1_a_ready;
	assign auto_tileClockGater_tile_clock_gater_in_d_valid = tileClockGater_auto_tile_clock_gater_in_1_d_valid;
	assign auto_tileClockGater_tile_clock_gater_in_d_bits_opcode = tileClockGater_auto_tile_clock_gater_in_1_d_bits_opcode;
	assign auto_tileClockGater_tile_clock_gater_in_d_bits_size = tileClockGater_auto_tile_clock_gater_in_1_d_bits_size;
	assign auto_tileClockGater_tile_clock_gater_in_d_bits_source = tileClockGater_auto_tile_clock_gater_in_1_d_bits_source;
	assign auto_tileClockGater_tile_clock_gater_in_d_bits_data = tileClockGater_auto_tile_clock_gater_in_1_d_bits_data;
	assign auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_clock = tileClockGater_auto_tile_clock_gater_out_member_allClocks_implicit_clock_clock;
	assign auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_reset = tileClockGater_auto_tile_clock_gater_out_member_allClocks_implicit_clock_reset;
	assign auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock = tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock;
	assign auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset = tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset;
	assign auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock = tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock;
	assign auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset = tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset;
	assign auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock = tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock;
	assign auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset = tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset;
	assign auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock = tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock;
	assign auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset = tileClockGater_auto_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset;
	assign tileClockGater_clock = auto_clock_in_clock;
	assign tileClockGater_reset = auto_clock_in_reset;
	assign tileClockGater_auto_tile_clock_gater_in_1_a_valid = auto_tileClockGater_tile_clock_gater_in_a_valid;
	assign tileClockGater_auto_tile_clock_gater_in_1_a_bits_opcode = auto_tileClockGater_tile_clock_gater_in_a_bits_opcode;
	assign tileClockGater_auto_tile_clock_gater_in_1_a_bits_param = auto_tileClockGater_tile_clock_gater_in_a_bits_param;
	assign tileClockGater_auto_tile_clock_gater_in_1_a_bits_size = auto_tileClockGater_tile_clock_gater_in_a_bits_size;
	assign tileClockGater_auto_tile_clock_gater_in_1_a_bits_source = auto_tileClockGater_tile_clock_gater_in_a_bits_source;
	assign tileClockGater_auto_tile_clock_gater_in_1_a_bits_address = auto_tileClockGater_tile_clock_gater_in_a_bits_address;
	assign tileClockGater_auto_tile_clock_gater_in_1_a_bits_mask = auto_tileClockGater_tile_clock_gater_in_a_bits_mask;
	assign tileClockGater_auto_tile_clock_gater_in_1_a_bits_data = auto_tileClockGater_tile_clock_gater_in_a_bits_data;
	assign tileClockGater_auto_tile_clock_gater_in_1_a_bits_corrupt = auto_tileClockGater_tile_clock_gater_in_a_bits_corrupt;
	assign tileClockGater_auto_tile_clock_gater_in_1_d_ready = auto_tileClockGater_tile_clock_gater_in_d_ready;
	assign tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_clock = tileResetSetter_auto_clock_out_member_allClocks_implicit_clock_clock;
	assign tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_implicit_clock_reset = tileResetSetter_auto_clock_out_member_allClocks_implicit_clock_reset;
	assign tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_clock = tileResetSetter_auto_clock_out_member_allClocks_subsystem_cbus_0_clock;
	assign tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_cbus_0_reset = tileResetSetter_auto_clock_out_member_allClocks_subsystem_cbus_0_reset;
	assign tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_clock = tileResetSetter_auto_clock_out_member_allClocks_subsystem_fbus_0_clock;
	assign tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_fbus_0_reset = tileResetSetter_auto_clock_out_member_allClocks_subsystem_fbus_0_reset;
	assign tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_clock = tileResetSetter_auto_clock_out_member_allClocks_subsystem_pbus_0_clock;
	assign tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_pbus_0_reset = tileResetSetter_auto_clock_out_member_allClocks_subsystem_pbus_0_reset;
	assign tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_clock = tileResetSetter_auto_clock_out_member_allClocks_subsystem_sbus_0_clock;
	assign tileClockGater_auto_tile_clock_gater_in_0_member_allClocks_subsystem_sbus_0_reset = tileResetSetter_auto_clock_out_member_allClocks_subsystem_sbus_0_reset;
	assign tileResetSetter_clock = auto_clock_in_clock;
	assign tileResetSetter_reset = auto_clock_in_reset;
	assign tileResetSetter_auto_clock_in_member_allClocks_implicit_clock_clock = auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock;
	assign tileResetSetter_auto_clock_in_member_allClocks_implicit_clock_reset = auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset;
	assign tileResetSetter_auto_clock_in_member_allClocks_subsystem_cbus_0_clock = auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock;
	assign tileResetSetter_auto_clock_in_member_allClocks_subsystem_cbus_0_reset = auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset;
	assign tileResetSetter_auto_clock_in_member_allClocks_subsystem_fbus_0_clock = auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock;
	assign tileResetSetter_auto_clock_in_member_allClocks_subsystem_fbus_0_reset = auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset;
	assign tileResetSetter_auto_clock_in_member_allClocks_subsystem_pbus_0_clock = auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock;
	assign tileResetSetter_auto_clock_in_member_allClocks_subsystem_pbus_0_reset = auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset;
	assign tileResetSetter_auto_clock_in_member_allClocks_subsystem_sbus_0_clock = auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock;
	assign tileResetSetter_auto_clock_in_member_allClocks_subsystem_sbus_0_reset = auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset;
	assign tileResetSetter_auto_tl_in_a_valid = auto_tileResetSetter_tl_in_a_valid;
	assign tileResetSetter_auto_tl_in_a_bits_opcode = auto_tileResetSetter_tl_in_a_bits_opcode;
	assign tileResetSetter_auto_tl_in_a_bits_param = auto_tileResetSetter_tl_in_a_bits_param;
	assign tileResetSetter_auto_tl_in_a_bits_size = auto_tileResetSetter_tl_in_a_bits_size;
	assign tileResetSetter_auto_tl_in_a_bits_source = auto_tileResetSetter_tl_in_a_bits_source;
	assign tileResetSetter_auto_tl_in_a_bits_address = auto_tileResetSetter_tl_in_a_bits_address;
	assign tileResetSetter_auto_tl_in_a_bits_mask = auto_tileResetSetter_tl_in_a_bits_mask;
	assign tileResetSetter_auto_tl_in_a_bits_data = auto_tileResetSetter_tl_in_a_bits_data;
	assign tileResetSetter_auto_tl_in_a_bits_corrupt = auto_tileResetSetter_tl_in_a_bits_corrupt;
	assign tileResetSetter_auto_tl_in_d_ready = auto_tileResetSetter_tl_in_d_ready;
endmodule
module ClockGroupAggregator_4 (
	auto_in_member_allClocks_implicit_clock_clock,
	auto_in_member_allClocks_implicit_clock_reset,
	auto_in_member_allClocks_subsystem_cbus_0_clock,
	auto_in_member_allClocks_subsystem_cbus_0_reset,
	auto_in_member_allClocks_subsystem_fbus_0_clock,
	auto_in_member_allClocks_subsystem_fbus_0_reset,
	auto_in_member_allClocks_subsystem_pbus_0_clock,
	auto_in_member_allClocks_subsystem_pbus_0_reset,
	auto_in_member_allClocks_subsystem_sbus_0_clock,
	auto_in_member_allClocks_subsystem_sbus_0_reset,
	auto_out_4_member_implicitClockGrouper_implicit_clock_clock,
	auto_out_4_member_implicitClockGrouper_implicit_clock_reset,
	auto_out_3_member_subsystem_cbus_subsystem_cbus_0_clock,
	auto_out_3_member_subsystem_cbus_subsystem_cbus_0_reset,
	auto_out_2_member_subsystem_fbus_subsystem_fbus_0_clock,
	auto_out_2_member_subsystem_fbus_subsystem_fbus_0_reset,
	auto_out_1_member_subsystem_pbus_subsystem_pbus_0_clock,
	auto_out_1_member_subsystem_pbus_subsystem_pbus_0_reset,
	auto_out_0_member_subsystem_sbus_subsystem_sbus_0_clock,
	auto_out_0_member_subsystem_sbus_subsystem_sbus_0_reset
);
	input auto_in_member_allClocks_implicit_clock_clock;
	input auto_in_member_allClocks_implicit_clock_reset;
	input auto_in_member_allClocks_subsystem_cbus_0_clock;
	input auto_in_member_allClocks_subsystem_cbus_0_reset;
	input auto_in_member_allClocks_subsystem_fbus_0_clock;
	input auto_in_member_allClocks_subsystem_fbus_0_reset;
	input auto_in_member_allClocks_subsystem_pbus_0_clock;
	input auto_in_member_allClocks_subsystem_pbus_0_reset;
	input auto_in_member_allClocks_subsystem_sbus_0_clock;
	input auto_in_member_allClocks_subsystem_sbus_0_reset;
	output wire auto_out_4_member_implicitClockGrouper_implicit_clock_clock;
	output wire auto_out_4_member_implicitClockGrouper_implicit_clock_reset;
	output wire auto_out_3_member_subsystem_cbus_subsystem_cbus_0_clock;
	output wire auto_out_3_member_subsystem_cbus_subsystem_cbus_0_reset;
	output wire auto_out_2_member_subsystem_fbus_subsystem_fbus_0_clock;
	output wire auto_out_2_member_subsystem_fbus_subsystem_fbus_0_reset;
	output wire auto_out_1_member_subsystem_pbus_subsystem_pbus_0_clock;
	output wire auto_out_1_member_subsystem_pbus_subsystem_pbus_0_reset;
	output wire auto_out_0_member_subsystem_sbus_subsystem_sbus_0_clock;
	output wire auto_out_0_member_subsystem_sbus_subsystem_sbus_0_reset;
	assign auto_out_4_member_implicitClockGrouper_implicit_clock_clock = auto_in_member_allClocks_implicit_clock_clock;
	assign auto_out_4_member_implicitClockGrouper_implicit_clock_reset = auto_in_member_allClocks_implicit_clock_reset;
	assign auto_out_3_member_subsystem_cbus_subsystem_cbus_0_clock = auto_in_member_allClocks_subsystem_cbus_0_clock;
	assign auto_out_3_member_subsystem_cbus_subsystem_cbus_0_reset = auto_in_member_allClocks_subsystem_cbus_0_reset;
	assign auto_out_2_member_subsystem_fbus_subsystem_fbus_0_clock = auto_in_member_allClocks_subsystem_fbus_0_clock;
	assign auto_out_2_member_subsystem_fbus_subsystem_fbus_0_reset = auto_in_member_allClocks_subsystem_fbus_0_reset;
	assign auto_out_1_member_subsystem_pbus_subsystem_pbus_0_clock = auto_in_member_allClocks_subsystem_pbus_0_clock;
	assign auto_out_1_member_subsystem_pbus_subsystem_pbus_0_reset = auto_in_member_allClocks_subsystem_pbus_0_reset;
	assign auto_out_0_member_subsystem_sbus_subsystem_sbus_0_clock = auto_in_member_allClocks_subsystem_sbus_0_clock;
	assign auto_out_0_member_subsystem_sbus_subsystem_sbus_0_reset = auto_in_member_allClocks_subsystem_sbus_0_reset;
endmodule
module ClockGroupParameterModifier (
	auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_clock,
	auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_reset,
	auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_clock,
	auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_reset,
	auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_clock,
	auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_reset,
	auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_clock,
	auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_reset,
	auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_clock,
	auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_reset,
	auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_clock,
	auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_reset,
	auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_clock,
	auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_reset,
	auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_clock,
	auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_reset
);
	input auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_clock;
	input auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_reset;
	input auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_clock;
	input auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_reset;
	input auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_clock;
	input auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_reset;
	input auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_clock;
	input auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_reset;
	output wire auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_clock;
	output wire auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_reset;
	output wire auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_clock;
	output wire auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_reset;
	output wire auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_clock;
	output wire auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_reset;
	output wire auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_clock;
	output wire auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_reset;
	assign auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_clock = auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_clock;
	assign auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_reset = auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_reset;
	assign auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_clock = auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_clock;
	assign auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_reset = auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_reset;
	assign auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_clock = auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_clock;
	assign auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_reset = auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_reset;
	assign auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_clock = auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_clock;
	assign auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_reset = auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_reset;
endmodule
module ClockGroupParameterModifier_1 (
	auto_frequency_specifier_in_member_allClocks_implicit_clock_clock,
	auto_frequency_specifier_in_member_allClocks_implicit_clock_reset,
	auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_clock,
	auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_reset,
	auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_clock,
	auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_reset,
	auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_clock,
	auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_reset,
	auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_clock,
	auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_reset,
	auto_frequency_specifier_out_member_allClocks_implicit_clock_clock,
	auto_frequency_specifier_out_member_allClocks_implicit_clock_reset,
	auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_clock,
	auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_reset,
	auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_clock,
	auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_reset,
	auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_clock,
	auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_reset,
	auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_clock,
	auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_reset
);
	input auto_frequency_specifier_in_member_allClocks_implicit_clock_clock;
	input auto_frequency_specifier_in_member_allClocks_implicit_clock_reset;
	input auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_clock;
	input auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_reset;
	input auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_clock;
	input auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_reset;
	input auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_clock;
	input auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_reset;
	input auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_clock;
	input auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_reset;
	output wire auto_frequency_specifier_out_member_allClocks_implicit_clock_clock;
	output wire auto_frequency_specifier_out_member_allClocks_implicit_clock_reset;
	output wire auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_clock;
	output wire auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_reset;
	output wire auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_clock;
	output wire auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_reset;
	output wire auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_clock;
	output wire auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_reset;
	output wire auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_clock;
	output wire auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_reset;
	assign auto_frequency_specifier_out_member_allClocks_implicit_clock_clock = auto_frequency_specifier_in_member_allClocks_implicit_clock_clock;
	assign auto_frequency_specifier_out_member_allClocks_implicit_clock_reset = auto_frequency_specifier_in_member_allClocks_implicit_clock_reset;
	assign auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_clock = auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_clock;
	assign auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_reset = auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_reset;
	assign auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_clock = auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_clock;
	assign auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_reset = auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_reset;
	assign auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_clock = auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_clock;
	assign auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_reset = auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_reset;
	assign auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_clock = auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_clock;
	assign auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_reset = auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_reset;
endmodule
module ClockGroupCombiner (
	auto_clock_group_combiner_in_member_allClocks_implicit_clock_clock,
	auto_clock_group_combiner_in_member_allClocks_implicit_clock_reset,
	auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_clock,
	auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_reset,
	auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_clock,
	auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_reset,
	auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_clock,
	auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_reset,
	auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_clock,
	auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_reset,
	auto_clock_group_combiner_out_member_allClocks_implicit_clock_clock,
	auto_clock_group_combiner_out_member_allClocks_implicit_clock_reset,
	auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_clock,
	auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_reset,
	auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_clock,
	auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_reset,
	auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_clock,
	auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_reset,
	auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_clock,
	auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_reset
);
	input auto_clock_group_combiner_in_member_allClocks_implicit_clock_clock;
	input auto_clock_group_combiner_in_member_allClocks_implicit_clock_reset;
	input auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_clock;
	input auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_reset;
	input auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_clock;
	input auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_reset;
	input auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_clock;
	input auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_reset;
	input auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_clock;
	input auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_reset;
	output wire auto_clock_group_combiner_out_member_allClocks_implicit_clock_clock;
	output wire auto_clock_group_combiner_out_member_allClocks_implicit_clock_reset;
	output wire auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_clock;
	output wire auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_reset;
	output wire auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_clock;
	output wire auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_reset;
	output wire auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_clock;
	output wire auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_reset;
	output wire auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_clock;
	output wire auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_reset;
	assign auto_clock_group_combiner_out_member_allClocks_implicit_clock_clock = auto_clock_group_combiner_in_member_allClocks_implicit_clock_clock;
	assign auto_clock_group_combiner_out_member_allClocks_implicit_clock_reset = auto_clock_group_combiner_in_member_allClocks_implicit_clock_reset;
	assign auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_clock = auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_clock;
	assign auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_reset = auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_reset;
	assign auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_clock = auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_clock;
	assign auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_reset = auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_reset;
	assign auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_clock = auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_clock;
	assign auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_reset = auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_reset;
	assign auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_clock = auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_clock;
	assign auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_reset = auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_reset;
endmodule
module ResetCatchAndSync_d3 (
	clock,
	reset,
	io_sync_reset
);
	input clock;
	input reset;
	output wire io_sync_reset;
	wire io_sync_reset_chain_clock;
	wire io_sync_reset_chain_reset;
	wire io_sync_reset_chain_io_d;
	wire io_sync_reset_chain_io_q;
	wire _io_sync_reset_WIRE = io_sync_reset_chain_io_q;
	AsyncResetSynchronizerShiftReg_w1_d3_i0 io_sync_reset_chain(
		.clock(io_sync_reset_chain_clock),
		.reset(io_sync_reset_chain_reset),
		.io_d(io_sync_reset_chain_io_d),
		.io_q(io_sync_reset_chain_io_q)
	);
	assign io_sync_reset = ~_io_sync_reset_WIRE;
	assign io_sync_reset_chain_clock = clock;
	assign io_sync_reset_chain_reset = reset;
	assign io_sync_reset_chain_io_d = 1'h1;
endmodule
module ClockGroupResetSynchronizer (
	auto_in_member_allClocks_implicit_clock_clock,
	auto_in_member_allClocks_implicit_clock_reset,
	auto_in_member_allClocks_subsystem_cbus_0_clock,
	auto_in_member_allClocks_subsystem_cbus_0_reset,
	auto_in_member_allClocks_subsystem_fbus_0_clock,
	auto_in_member_allClocks_subsystem_fbus_0_reset,
	auto_in_member_allClocks_subsystem_pbus_0_clock,
	auto_in_member_allClocks_subsystem_pbus_0_reset,
	auto_in_member_allClocks_subsystem_sbus_0_clock,
	auto_in_member_allClocks_subsystem_sbus_0_reset,
	auto_out_member_allClocks_implicit_clock_clock,
	auto_out_member_allClocks_implicit_clock_reset,
	auto_out_member_allClocks_subsystem_cbus_0_clock,
	auto_out_member_allClocks_subsystem_cbus_0_reset,
	auto_out_member_allClocks_subsystem_fbus_0_clock,
	auto_out_member_allClocks_subsystem_fbus_0_reset,
	auto_out_member_allClocks_subsystem_pbus_0_clock,
	auto_out_member_allClocks_subsystem_pbus_0_reset,
	auto_out_member_allClocks_subsystem_sbus_0_clock,
	auto_out_member_allClocks_subsystem_sbus_0_reset
);
	input auto_in_member_allClocks_implicit_clock_clock;
	input auto_in_member_allClocks_implicit_clock_reset;
	input auto_in_member_allClocks_subsystem_cbus_0_clock;
	input auto_in_member_allClocks_subsystem_cbus_0_reset;
	input auto_in_member_allClocks_subsystem_fbus_0_clock;
	input auto_in_member_allClocks_subsystem_fbus_0_reset;
	input auto_in_member_allClocks_subsystem_pbus_0_clock;
	input auto_in_member_allClocks_subsystem_pbus_0_reset;
	input auto_in_member_allClocks_subsystem_sbus_0_clock;
	input auto_in_member_allClocks_subsystem_sbus_0_reset;
	output wire auto_out_member_allClocks_implicit_clock_clock;
	output wire auto_out_member_allClocks_implicit_clock_reset;
	output wire auto_out_member_allClocks_subsystem_cbus_0_clock;
	output wire auto_out_member_allClocks_subsystem_cbus_0_reset;
	output wire auto_out_member_allClocks_subsystem_fbus_0_clock;
	output wire auto_out_member_allClocks_subsystem_fbus_0_reset;
	output wire auto_out_member_allClocks_subsystem_pbus_0_clock;
	output wire auto_out_member_allClocks_subsystem_pbus_0_reset;
	output wire auto_out_member_allClocks_subsystem_sbus_0_clock;
	output wire auto_out_member_allClocks_subsystem_sbus_0_reset;
	wire bundleOut_0_member_allClocks_subsystem_sbus_0_reset_catcher_clock;
	wire bundleOut_0_member_allClocks_subsystem_sbus_0_reset_catcher_reset;
	wire bundleOut_0_member_allClocks_subsystem_sbus_0_reset_catcher_io_sync_reset;
	wire bundleOut_0_member_allClocks_subsystem_pbus_0_reset_catcher_clock;
	wire bundleOut_0_member_allClocks_subsystem_pbus_0_reset_catcher_reset;
	wire bundleOut_0_member_allClocks_subsystem_pbus_0_reset_catcher_io_sync_reset;
	wire bundleOut_0_member_allClocks_subsystem_fbus_0_reset_catcher_clock;
	wire bundleOut_0_member_allClocks_subsystem_fbus_0_reset_catcher_reset;
	wire bundleOut_0_member_allClocks_subsystem_fbus_0_reset_catcher_io_sync_reset;
	wire bundleOut_0_member_allClocks_subsystem_cbus_0_reset_catcher_clock;
	wire bundleOut_0_member_allClocks_subsystem_cbus_0_reset_catcher_reset;
	wire bundleOut_0_member_allClocks_subsystem_cbus_0_reset_catcher_io_sync_reset;
	wire bundleOut_0_member_allClocks_implicit_clock_reset_catcher_clock;
	wire bundleOut_0_member_allClocks_implicit_clock_reset_catcher_reset;
	wire bundleOut_0_member_allClocks_implicit_clock_reset_catcher_io_sync_reset;
	ResetCatchAndSync_d3 bundleOut_0_member_allClocks_subsystem_sbus_0_reset_catcher(
		.clock(bundleOut_0_member_allClocks_subsystem_sbus_0_reset_catcher_clock),
		.reset(bundleOut_0_member_allClocks_subsystem_sbus_0_reset_catcher_reset),
		.io_sync_reset(bundleOut_0_member_allClocks_subsystem_sbus_0_reset_catcher_io_sync_reset)
	);
	ResetCatchAndSync_d3 bundleOut_0_member_allClocks_subsystem_pbus_0_reset_catcher(
		.clock(bundleOut_0_member_allClocks_subsystem_pbus_0_reset_catcher_clock),
		.reset(bundleOut_0_member_allClocks_subsystem_pbus_0_reset_catcher_reset),
		.io_sync_reset(bundleOut_0_member_allClocks_subsystem_pbus_0_reset_catcher_io_sync_reset)
	);
	ResetCatchAndSync_d3 bundleOut_0_member_allClocks_subsystem_fbus_0_reset_catcher(
		.clock(bundleOut_0_member_allClocks_subsystem_fbus_0_reset_catcher_clock),
		.reset(bundleOut_0_member_allClocks_subsystem_fbus_0_reset_catcher_reset),
		.io_sync_reset(bundleOut_0_member_allClocks_subsystem_fbus_0_reset_catcher_io_sync_reset)
	);
	ResetCatchAndSync_d3 bundleOut_0_member_allClocks_subsystem_cbus_0_reset_catcher(
		.clock(bundleOut_0_member_allClocks_subsystem_cbus_0_reset_catcher_clock),
		.reset(bundleOut_0_member_allClocks_subsystem_cbus_0_reset_catcher_reset),
		.io_sync_reset(bundleOut_0_member_allClocks_subsystem_cbus_0_reset_catcher_io_sync_reset)
	);
	ResetCatchAndSync_d3 bundleOut_0_member_allClocks_implicit_clock_reset_catcher(
		.clock(bundleOut_0_member_allClocks_implicit_clock_reset_catcher_clock),
		.reset(bundleOut_0_member_allClocks_implicit_clock_reset_catcher_reset),
		.io_sync_reset(bundleOut_0_member_allClocks_implicit_clock_reset_catcher_io_sync_reset)
	);
	assign auto_out_member_allClocks_implicit_clock_clock = auto_in_member_allClocks_implicit_clock_clock;
	assign auto_out_member_allClocks_implicit_clock_reset = bundleOut_0_member_allClocks_implicit_clock_reset_catcher_io_sync_reset;
	assign auto_out_member_allClocks_subsystem_cbus_0_clock = auto_in_member_allClocks_subsystem_cbus_0_clock;
	assign auto_out_member_allClocks_subsystem_cbus_0_reset = bundleOut_0_member_allClocks_subsystem_cbus_0_reset_catcher_io_sync_reset;
	assign auto_out_member_allClocks_subsystem_fbus_0_clock = auto_in_member_allClocks_subsystem_fbus_0_clock;
	assign auto_out_member_allClocks_subsystem_fbus_0_reset = bundleOut_0_member_allClocks_subsystem_fbus_0_reset_catcher_io_sync_reset;
	assign auto_out_member_allClocks_subsystem_pbus_0_clock = auto_in_member_allClocks_subsystem_pbus_0_clock;
	assign auto_out_member_allClocks_subsystem_pbus_0_reset = bundleOut_0_member_allClocks_subsystem_pbus_0_reset_catcher_io_sync_reset;
	assign auto_out_member_allClocks_subsystem_sbus_0_clock = auto_in_member_allClocks_subsystem_sbus_0_clock;
	assign auto_out_member_allClocks_subsystem_sbus_0_reset = bundleOut_0_member_allClocks_subsystem_sbus_0_reset_catcher_io_sync_reset;
	assign bundleOut_0_member_allClocks_subsystem_sbus_0_reset_catcher_clock = auto_in_member_allClocks_subsystem_sbus_0_clock;
	assign bundleOut_0_member_allClocks_subsystem_sbus_0_reset_catcher_reset = auto_in_member_allClocks_subsystem_sbus_0_reset;
	assign bundleOut_0_member_allClocks_subsystem_pbus_0_reset_catcher_clock = auto_in_member_allClocks_subsystem_pbus_0_clock;
	assign bundleOut_0_member_allClocks_subsystem_pbus_0_reset_catcher_reset = auto_in_member_allClocks_subsystem_pbus_0_reset;
	assign bundleOut_0_member_allClocks_subsystem_fbus_0_reset_catcher_clock = auto_in_member_allClocks_subsystem_fbus_0_clock;
	assign bundleOut_0_member_allClocks_subsystem_fbus_0_reset_catcher_reset = auto_in_member_allClocks_subsystem_fbus_0_reset;
	assign bundleOut_0_member_allClocks_subsystem_cbus_0_reset_catcher_clock = auto_in_member_allClocks_subsystem_cbus_0_clock;
	assign bundleOut_0_member_allClocks_subsystem_cbus_0_reset_catcher_reset = auto_in_member_allClocks_subsystem_cbus_0_reset;
	assign bundleOut_0_member_allClocks_implicit_clock_reset_catcher_clock = auto_in_member_allClocks_implicit_clock_clock;
	assign bundleOut_0_member_allClocks_implicit_clock_reset_catcher_reset = auto_in_member_allClocks_implicit_clock_reset;
endmodule
module ClockGroup_4 (
	auto_in_member_implicitClockGrouper_implicit_clock_clock,
	auto_in_member_implicitClockGrouper_implicit_clock_reset,
	auto_out_clock,
	auto_out_reset
);
	input auto_in_member_implicitClockGrouper_implicit_clock_clock;
	input auto_in_member_implicitClockGrouper_implicit_clock_reset;
	output wire auto_out_clock;
	output wire auto_out_reset;
	assign auto_out_clock = auto_in_member_implicitClockGrouper_implicit_clock_clock;
	assign auto_out_reset = auto_in_member_implicitClockGrouper_implicit_clock_reset;
endmodule
module CaptureUpdateChain (
	clock,
	reset,
	io_chainIn_shift,
	io_chainIn_data,
	io_chainIn_capture,
	io_chainIn_update,
	io_chainOut_data,
	io_capture_bits_dmiStatus,
	io_update_valid,
	io_update_bits_dmireset
);
	input clock;
	input reset;
	input io_chainIn_shift;
	input io_chainIn_data;
	input io_chainIn_capture;
	input io_chainIn_update;
	output wire io_chainOut_data;
	input [1:0] io_capture_bits_dmiStatus;
	output wire io_update_valid;
	output wire io_update_bits_dmireset;
	reg regs_0;
	reg regs_1;
	reg regs_2;
	reg regs_3;
	reg regs_4;
	reg regs_5;
	reg regs_6;
	reg regs_7;
	reg regs_8;
	reg regs_9;
	reg regs_10;
	reg regs_11;
	reg regs_12;
	reg regs_13;
	reg regs_14;
	reg regs_15;
	reg regs_16;
	reg regs_17;
	reg regs_18;
	reg regs_19;
	reg regs_20;
	reg regs_21;
	reg regs_22;
	reg regs_23;
	reg regs_24;
	reg regs_25;
	reg regs_26;
	reg regs_27;
	reg regs_28;
	reg regs_29;
	reg regs_30;
	reg regs_31;
	wire [7:0] updateBits_lo_lo = {regs_7, regs_6, regs_5, regs_4, regs_3, regs_2, regs_1, regs_0};
	wire [15:0] updateBits_lo = {regs_15, regs_14, regs_13, regs_12, regs_11, regs_10, regs_9, regs_8, updateBits_lo_lo};
	wire [7:0] updateBits_hi_lo = {regs_23, regs_22, regs_21, regs_20, regs_19, regs_18, regs_17, regs_16};
	wire [31:0] updateBits = {regs_31, regs_30, regs_29, regs_28, regs_27, regs_26, regs_25, regs_24, updateBits_hi_lo, updateBits_lo};
	wire [31:0] captureBits = {20'h00005, io_capture_bits_dmiStatus, 6'h07, 4'h1};
	wire _T_1 = ~(io_chainIn_capture & io_chainIn_update);
	wire _T_4 = _T_1 & ~(io_chainIn_capture & io_chainIn_shift);
	wire _T_7 = _T_4 & ~(io_chainIn_update & io_chainIn_shift);
	assign io_chainOut_data = regs_0;
	assign io_update_valid = (io_chainIn_capture ? 1'h0 : io_chainIn_update);
	assign io_update_bits_dmireset = updateBits[16];
	always @(posedge clock) begin
		if (io_chainIn_capture)
			regs_0 <= captureBits[0];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_0 <= regs_1;
		if (io_chainIn_capture)
			regs_1 <= captureBits[1];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_1 <= regs_2;
		if (io_chainIn_capture)
			regs_2 <= captureBits[2];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_2 <= regs_3;
		if (io_chainIn_capture)
			regs_3 <= captureBits[3];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_3 <= regs_4;
		if (io_chainIn_capture)
			regs_4 <= captureBits[4];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_4 <= regs_5;
		if (io_chainIn_capture)
			regs_5 <= captureBits[5];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_5 <= regs_6;
		if (io_chainIn_capture)
			regs_6 <= captureBits[6];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_6 <= regs_7;
		if (io_chainIn_capture)
			regs_7 <= captureBits[7];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_7 <= regs_8;
		if (io_chainIn_capture)
			regs_8 <= captureBits[8];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_8 <= regs_9;
		if (io_chainIn_capture)
			regs_9 <= captureBits[9];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_9 <= regs_10;
		if (io_chainIn_capture)
			regs_10 <= captureBits[10];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_10 <= regs_11;
		if (io_chainIn_capture)
			regs_11 <= captureBits[11];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_11 <= regs_12;
		if (io_chainIn_capture)
			regs_12 <= captureBits[12];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_12 <= regs_13;
		if (io_chainIn_capture)
			regs_13 <= captureBits[13];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_13 <= regs_14;
		if (io_chainIn_capture)
			regs_14 <= captureBits[14];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_14 <= regs_15;
		if (io_chainIn_capture)
			regs_15 <= captureBits[15];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_15 <= regs_16;
		if (io_chainIn_capture)
			regs_16 <= captureBits[16];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_16 <= regs_17;
		if (io_chainIn_capture)
			regs_17 <= captureBits[17];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_17 <= regs_18;
		if (io_chainIn_capture)
			regs_18 <= captureBits[18];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_18 <= regs_19;
		if (io_chainIn_capture)
			regs_19 <= captureBits[19];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_19 <= regs_20;
		if (io_chainIn_capture)
			regs_20 <= captureBits[20];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_20 <= regs_21;
		if (io_chainIn_capture)
			regs_21 <= captureBits[21];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_21 <= regs_22;
		if (io_chainIn_capture)
			regs_22 <= captureBits[22];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_22 <= regs_23;
		if (io_chainIn_capture)
			regs_23 <= captureBits[23];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_23 <= regs_24;
		if (io_chainIn_capture)
			regs_24 <= captureBits[24];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_24 <= regs_25;
		if (io_chainIn_capture)
			regs_25 <= captureBits[25];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_25 <= regs_26;
		if (io_chainIn_capture)
			regs_26 <= captureBits[26];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_26 <= regs_27;
		if (io_chainIn_capture)
			regs_27 <= captureBits[27];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_27 <= regs_28;
		if (io_chainIn_capture)
			regs_28 <= captureBits[28];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_28 <= regs_29;
		if (io_chainIn_capture)
			regs_29 <= captureBits[29];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_29 <= regs_30;
		if (io_chainIn_capture)
			regs_30 <= captureBits[30];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_30 <= regs_31;
		if (io_chainIn_capture)
			regs_31 <= captureBits[31];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_31 <= io_chainIn_data;
	end
endmodule
module CaptureUpdateChain_1 (
	clock,
	reset,
	io_chainIn_shift,
	io_chainIn_data,
	io_chainIn_capture,
	io_chainIn_update,
	io_chainOut_data,
	io_capture_bits_addr,
	io_capture_bits_data,
	io_capture_bits_resp,
	io_capture_capture,
	io_update_valid,
	io_update_bits_addr,
	io_update_bits_data,
	io_update_bits_op
);
	input clock;
	input reset;
	input io_chainIn_shift;
	input io_chainIn_data;
	input io_chainIn_capture;
	input io_chainIn_update;
	output wire io_chainOut_data;
	input [6:0] io_capture_bits_addr;
	input [31:0] io_capture_bits_data;
	input [1:0] io_capture_bits_resp;
	output wire io_capture_capture;
	output wire io_update_valid;
	output wire [6:0] io_update_bits_addr;
	output wire [31:0] io_update_bits_data;
	output wire [1:0] io_update_bits_op;
	reg regs_0;
	reg regs_1;
	reg regs_2;
	reg regs_3;
	reg regs_4;
	reg regs_5;
	reg regs_6;
	reg regs_7;
	reg regs_8;
	reg regs_9;
	reg regs_10;
	reg regs_11;
	reg regs_12;
	reg regs_13;
	reg regs_14;
	reg regs_15;
	reg regs_16;
	reg regs_17;
	reg regs_18;
	reg regs_19;
	reg regs_20;
	reg regs_21;
	reg regs_22;
	reg regs_23;
	reg regs_24;
	reg regs_25;
	reg regs_26;
	reg regs_27;
	reg regs_28;
	reg regs_29;
	reg regs_30;
	reg regs_31;
	reg regs_32;
	reg regs_33;
	reg regs_34;
	reg regs_35;
	reg regs_36;
	reg regs_37;
	reg regs_38;
	reg regs_39;
	reg regs_40;
	wire [9:0] updateBits_lo_lo = {regs_9, regs_8, regs_7, regs_6, regs_5, regs_4, regs_3, regs_2, regs_1, regs_0};
	wire [9:0] updateBits_lo_hi = {regs_19, regs_18, regs_17, regs_16, regs_15, regs_14, regs_13, regs_12, regs_11, regs_10};
	wire [9:0] updateBits_hi_lo = {regs_29, regs_28, regs_27, regs_26, regs_25, regs_24, regs_23, regs_22, regs_21, regs_20};
	wire [4:0] updateBits_hi_hi_lo = {regs_34, regs_33, regs_32, regs_31, regs_30};
	wire [40:0] updateBits = {regs_40, regs_39, regs_38, regs_37, regs_36, regs_35, updateBits_hi_hi_lo, updateBits_hi_lo, updateBits_lo_hi, updateBits_lo_lo};
	wire [40:0] captureBits = {io_capture_bits_addr, io_capture_bits_data, io_capture_bits_resp};
	wire _T_1 = ~(io_chainIn_capture & io_chainIn_update);
	wire _T_4 = _T_1 & ~(io_chainIn_capture & io_chainIn_shift);
	wire _T_7 = _T_4 & ~(io_chainIn_update & io_chainIn_shift);
	assign io_chainOut_data = regs_0;
	assign io_capture_capture = io_chainIn_capture;
	assign io_update_valid = (io_chainIn_capture ? 1'h0 : io_chainIn_update);
	assign io_update_bits_addr = updateBits[40:34];
	assign io_update_bits_data = updateBits[33:2];
	assign io_update_bits_op = updateBits[1:0];
	always @(posedge clock) begin
		if (io_chainIn_capture)
			regs_0 <= captureBits[0];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_0 <= regs_1;
		if (io_chainIn_capture)
			regs_1 <= captureBits[1];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_1 <= regs_2;
		if (io_chainIn_capture)
			regs_2 <= captureBits[2];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_2 <= regs_3;
		if (io_chainIn_capture)
			regs_3 <= captureBits[3];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_3 <= regs_4;
		if (io_chainIn_capture)
			regs_4 <= captureBits[4];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_4 <= regs_5;
		if (io_chainIn_capture)
			regs_5 <= captureBits[5];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_5 <= regs_6;
		if (io_chainIn_capture)
			regs_6 <= captureBits[6];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_6 <= regs_7;
		if (io_chainIn_capture)
			regs_7 <= captureBits[7];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_7 <= regs_8;
		if (io_chainIn_capture)
			regs_8 <= captureBits[8];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_8 <= regs_9;
		if (io_chainIn_capture)
			regs_9 <= captureBits[9];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_9 <= regs_10;
		if (io_chainIn_capture)
			regs_10 <= captureBits[10];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_10 <= regs_11;
		if (io_chainIn_capture)
			regs_11 <= captureBits[11];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_11 <= regs_12;
		if (io_chainIn_capture)
			regs_12 <= captureBits[12];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_12 <= regs_13;
		if (io_chainIn_capture)
			regs_13 <= captureBits[13];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_13 <= regs_14;
		if (io_chainIn_capture)
			regs_14 <= captureBits[14];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_14 <= regs_15;
		if (io_chainIn_capture)
			regs_15 <= captureBits[15];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_15 <= regs_16;
		if (io_chainIn_capture)
			regs_16 <= captureBits[16];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_16 <= regs_17;
		if (io_chainIn_capture)
			regs_17 <= captureBits[17];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_17 <= regs_18;
		if (io_chainIn_capture)
			regs_18 <= captureBits[18];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_18 <= regs_19;
		if (io_chainIn_capture)
			regs_19 <= captureBits[19];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_19 <= regs_20;
		if (io_chainIn_capture)
			regs_20 <= captureBits[20];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_20 <= regs_21;
		if (io_chainIn_capture)
			regs_21 <= captureBits[21];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_21 <= regs_22;
		if (io_chainIn_capture)
			regs_22 <= captureBits[22];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_22 <= regs_23;
		if (io_chainIn_capture)
			regs_23 <= captureBits[23];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_23 <= regs_24;
		if (io_chainIn_capture)
			regs_24 <= captureBits[24];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_24 <= regs_25;
		if (io_chainIn_capture)
			regs_25 <= captureBits[25];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_25 <= regs_26;
		if (io_chainIn_capture)
			regs_26 <= captureBits[26];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_26 <= regs_27;
		if (io_chainIn_capture)
			regs_27 <= captureBits[27];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_27 <= regs_28;
		if (io_chainIn_capture)
			regs_28 <= captureBits[28];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_28 <= regs_29;
		if (io_chainIn_capture)
			regs_29 <= captureBits[29];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_29 <= regs_30;
		if (io_chainIn_capture)
			regs_30 <= captureBits[30];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_30 <= regs_31;
		if (io_chainIn_capture)
			regs_31 <= captureBits[31];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_31 <= regs_32;
		if (io_chainIn_capture)
			regs_32 <= captureBits[32];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_32 <= regs_33;
		if (io_chainIn_capture)
			regs_33 <= captureBits[33];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_33 <= regs_34;
		if (io_chainIn_capture)
			regs_34 <= captureBits[34];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_34 <= regs_35;
		if (io_chainIn_capture)
			regs_35 <= captureBits[35];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_35 <= regs_36;
		if (io_chainIn_capture)
			regs_36 <= captureBits[36];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_36 <= regs_37;
		if (io_chainIn_capture)
			regs_37 <= captureBits[37];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_37 <= regs_38;
		if (io_chainIn_capture)
			regs_38 <= captureBits[38];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_38 <= regs_39;
		if (io_chainIn_capture)
			regs_39 <= captureBits[39];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_39 <= regs_40;
		if (io_chainIn_capture)
			regs_40 <= captureBits[40];
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_40 <= io_chainIn_data;
	end
endmodule
module CaptureChain (
	clock,
	reset,
	io_chainIn_shift,
	io_chainIn_data,
	io_chainIn_capture,
	io_chainIn_update,
	io_chainOut_data
);
	input clock;
	input reset;
	input io_chainIn_shift;
	input io_chainIn_data;
	input io_chainIn_capture;
	input io_chainIn_update;
	output wire io_chainOut_data;
	reg regs_0;
	reg regs_1;
	reg regs_2;
	reg regs_3;
	reg regs_4;
	reg regs_5;
	reg regs_6;
	reg regs_7;
	reg regs_8;
	reg regs_9;
	reg regs_10;
	reg regs_11;
	reg regs_12;
	reg regs_13;
	reg regs_14;
	reg regs_15;
	reg regs_16;
	reg regs_17;
	reg regs_18;
	reg regs_19;
	reg regs_20;
	reg regs_21;
	reg regs_22;
	reg regs_23;
	reg regs_24;
	reg regs_25;
	reg regs_26;
	reg regs_27;
	reg regs_28;
	reg regs_29;
	reg regs_30;
	reg regs_31;
	wire _GEN_1 = (io_chainIn_shift ? regs_1 : regs_0);
	wire _T_1 = ~(io_chainIn_capture & io_chainIn_update);
	wire _T_4 = _T_1 & ~(io_chainIn_capture & io_chainIn_shift);
	wire _T_7 = _T_4 & ~(io_chainIn_update & io_chainIn_shift);
	assign io_chainOut_data = regs_0;
	always @(posedge clock) begin
		regs_0 <= io_chainIn_capture | _GEN_1;
		if (io_chainIn_capture)
			regs_1 <= 1'h0;
		else if (io_chainIn_shift)
			regs_1 <= regs_2;
		if (io_chainIn_capture)
			regs_2 <= 1'h0;
		else if (io_chainIn_shift)
			regs_2 <= regs_3;
		if (io_chainIn_capture)
			regs_3 <= 1'h0;
		else if (io_chainIn_shift)
			regs_3 <= regs_4;
		if (io_chainIn_capture)
			regs_4 <= 1'h0;
		else if (io_chainIn_shift)
			regs_4 <= regs_5;
		if (io_chainIn_capture)
			regs_5 <= 1'h0;
		else if (io_chainIn_shift)
			regs_5 <= regs_6;
		if (io_chainIn_capture)
			regs_6 <= 1'h0;
		else if (io_chainIn_shift)
			regs_6 <= regs_7;
		if (io_chainIn_capture)
			regs_7 <= 1'h0;
		else if (io_chainIn_shift)
			regs_7 <= regs_8;
		if (io_chainIn_capture)
			regs_8 <= 1'h0;
		else if (io_chainIn_shift)
			regs_8 <= regs_9;
		if (io_chainIn_capture)
			regs_9 <= 1'h0;
		else if (io_chainIn_shift)
			regs_9 <= regs_10;
		if (io_chainIn_capture)
			regs_10 <= 1'h0;
		else if (io_chainIn_shift)
			regs_10 <= regs_11;
		if (io_chainIn_capture)
			regs_11 <= 1'h0;
		else if (io_chainIn_shift)
			regs_11 <= regs_12;
		if (io_chainIn_capture)
			regs_12 <= 1'h0;
		else if (io_chainIn_shift)
			regs_12 <= regs_13;
		if (io_chainIn_capture)
			regs_13 <= 1'h0;
		else if (io_chainIn_shift)
			regs_13 <= regs_14;
		if (io_chainIn_capture)
			regs_14 <= 1'h0;
		else if (io_chainIn_shift)
			regs_14 <= regs_15;
		if (io_chainIn_capture)
			regs_15 <= 1'h0;
		else if (io_chainIn_shift)
			regs_15 <= regs_16;
		if (io_chainIn_capture)
			regs_16 <= 1'h0;
		else if (io_chainIn_shift)
			regs_16 <= regs_17;
		if (io_chainIn_capture)
			regs_17 <= 1'h0;
		else if (io_chainIn_shift)
			regs_17 <= regs_18;
		if (io_chainIn_capture)
			regs_18 <= 1'h0;
		else if (io_chainIn_shift)
			regs_18 <= regs_19;
		if (io_chainIn_capture)
			regs_19 <= 1'h0;
		else if (io_chainIn_shift)
			regs_19 <= regs_20;
		if (io_chainIn_capture)
			regs_20 <= 1'h0;
		else if (io_chainIn_shift)
			regs_20 <= regs_21;
		if (io_chainIn_capture)
			regs_21 <= 1'h0;
		else if (io_chainIn_shift)
			regs_21 <= regs_22;
		if (io_chainIn_capture)
			regs_22 <= 1'h0;
		else if (io_chainIn_shift)
			regs_22 <= regs_23;
		if (io_chainIn_capture)
			regs_23 <= 1'h0;
		else if (io_chainIn_shift)
			regs_23 <= regs_24;
		if (io_chainIn_capture)
			regs_24 <= 1'h0;
		else if (io_chainIn_shift)
			regs_24 <= regs_25;
		if (io_chainIn_capture)
			regs_25 <= 1'h0;
		else if (io_chainIn_shift)
			regs_25 <= regs_26;
		if (io_chainIn_capture)
			regs_26 <= 1'h0;
		else if (io_chainIn_shift)
			regs_26 <= regs_27;
		if (io_chainIn_capture)
			regs_27 <= 1'h0;
		else if (io_chainIn_shift)
			regs_27 <= regs_28;
		if (io_chainIn_capture)
			regs_28 <= 1'h0;
		else if (io_chainIn_shift)
			regs_28 <= regs_29;
		if (io_chainIn_capture)
			regs_29 <= 1'h0;
		else if (io_chainIn_shift)
			regs_29 <= regs_30;
		if (io_chainIn_capture)
			regs_30 <= 1'h0;
		else if (io_chainIn_shift)
			regs_30 <= regs_31;
		if (io_chainIn_capture)
			regs_31 <= 1'h0;
		else if (io_chainIn_shift)
			regs_31 <= io_chainIn_data;
	end
endmodule
module JtagStateMachine (
	clock,
	reset,
	io_tms,
	io_currState
);
	input clock;
	input reset;
	input io_tms;
	output wire [3:0] io_currState;
	reg [3:0] currState;
	wire [3:0] _nextState_T_1 = (io_tms ? 4'h7 : 4'hc);
	wire [3:0] _nextState_T_3 = (io_tms ? 4'h1 : 4'h2);
	wire [3:0] _nextState_T_5 = (io_tms ? 4'h5 : 4'h3);
	wire [3:0] _nextState_T_6 = (io_tms ? 4'h0 : 4'h3);
	wire [3:0] _nextState_T_7 = (io_tms ? 4'h5 : 4'h2);
	wire [3:0] _nextState_T_9 = (io_tms ? 4'hf : 4'he);
	wire [3:0] _nextState_T_10 = (io_tms ? 4'h9 : 4'ha);
	wire [3:0] _nextState_T_12 = (io_tms ? 4'hd : 4'hb);
	wire [3:0] _nextState_T_13 = (io_tms ? 4'h8 : 4'hb);
	wire [3:0] _nextState_T_14 = (io_tms ? 4'hd : 4'ha);
	wire [3:0] _GEN_0 = (4'hd == currState ? _nextState_T_1 : 4'hf);
	wire [3:0] _GEN_1 = (4'h8 == currState ? _nextState_T_14 : _GEN_0);
	wire [3:0] _GEN_2 = (4'hb == currState ? _nextState_T_13 : _GEN_1);
	wire [3:0] _GEN_3 = (4'h9 == currState ? _nextState_T_12 : _GEN_2);
	wire [3:0] _GEN_4 = (4'ha == currState ? _nextState_T_10 : _GEN_3);
	wire [3:0] _GEN_5 = (4'he == currState ? _nextState_T_10 : _GEN_4);
	wire [3:0] _GEN_6 = (4'h4 == currState ? _nextState_T_9 : _GEN_5);
	wire [3:0] _GEN_7 = (4'h5 == currState ? _nextState_T_1 : _GEN_6);
	wire [3:0] _GEN_8 = (4'h0 == currState ? _nextState_T_7 : _GEN_7);
	wire [3:0] _GEN_9 = (4'h3 == currState ? _nextState_T_6 : _GEN_8);
	wire [3:0] _GEN_10 = (4'h1 == currState ? _nextState_T_5 : _GEN_9);
	wire [3:0] _GEN_11 = (4'h2 == currState ? _nextState_T_3 : _GEN_10);
	assign io_currState = currState;
	always @(posedge clock or posedge reset)
		if (reset)
			currState <= 4'hf;
		else if (4'hf == currState) begin
			if (io_tms)
				currState <= 4'hf;
			else
				currState <= 4'hc;
		end
		else if (4'hc == currState) begin
			if (io_tms)
				currState <= 4'h7;
			else
				currState <= 4'hc;
		end
		else if (4'h7 == currState) begin
			if (io_tms)
				currState <= 4'h4;
			else
				currState <= 4'h6;
		end
		else if (4'h6 == currState)
			currState <= _nextState_T_3;
		else
			currState <= _GEN_11;
endmodule
module CaptureUpdateChain_2 (
	clock,
	reset,
	io_chainIn_shift,
	io_chainIn_data,
	io_chainIn_capture,
	io_chainIn_update,
	io_chainOut_data,
	io_update_bits
);
	input clock;
	input reset;
	input io_chainIn_shift;
	input io_chainIn_data;
	input io_chainIn_capture;
	input io_chainIn_update;
	output wire io_chainOut_data;
	output wire [4:0] io_update_bits;
	reg regs_0;
	reg regs_1;
	reg regs_2;
	reg regs_3;
	reg regs_4;
	wire [1:0] updateBits_lo = {regs_1, regs_0};
	wire [2:0] updateBits_hi = {regs_4, regs_3, regs_2};
	wire _GEN_1 = (io_chainIn_shift ? regs_1 : regs_0);
	wire _GEN_9 = (io_chainIn_update ? regs_0 : _GEN_1);
	wire _T_1 = ~(io_chainIn_capture & io_chainIn_update);
	wire _T_4 = _T_1 & ~(io_chainIn_capture & io_chainIn_shift);
	wire _T_7 = _T_4 & ~(io_chainIn_update & io_chainIn_shift);
	assign io_chainOut_data = regs_0;
	assign io_update_bits = {updateBits_hi, updateBits_lo};
	always @(posedge clock) begin
		regs_0 <= io_chainIn_capture | _GEN_9;
		if (io_chainIn_capture)
			regs_1 <= 1'h0;
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_1 <= regs_2;
		if (io_chainIn_capture)
			regs_2 <= 1'h0;
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_2 <= regs_3;
		if (io_chainIn_capture)
			regs_3 <= 1'h0;
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_3 <= regs_4;
		if (io_chainIn_capture)
			regs_4 <= 1'h0;
		else if (!io_chainIn_update)
			if (io_chainIn_shift)
				regs_4 <= io_chainIn_data;
	end
endmodule
module JtagTapController (
	clock,
	reset,
	io_jtag_TMS,
	io_jtag_TDI,
	io_jtag_TDO_data,
	io_control_jtag_reset,
	io_output_instruction,
	io_output_tapIsInTestLogicReset,
	io_dataChainOut_shift,
	io_dataChainOut_data,
	io_dataChainOut_capture,
	io_dataChainOut_update,
	io_dataChainIn_data
);
	input clock;
	input reset;
	input io_jtag_TMS;
	input io_jtag_TDI;
	output wire io_jtag_TDO_data;
	input io_control_jtag_reset;
	output wire [4:0] io_output_instruction;
	output wire io_output_tapIsInTestLogicReset;
	output wire io_dataChainOut_shift;
	output wire io_dataChainOut_data;
	output wire io_dataChainOut_capture;
	output wire io_dataChainOut_update;
	input io_dataChainIn_data;
	wire stateMachine_clock;
	wire stateMachine_reset;
	wire stateMachine_io_tms;
	wire [3:0] stateMachine_io_currState;
	wire irChain_clock;
	wire irChain_reset;
	wire irChain_io_chainIn_shift;
	wire irChain_io_chainIn_data;
	wire irChain_io_chainIn_capture;
	wire irChain_io_chainIn_update;
	wire irChain_io_chainOut_data;
	wire [4:0] irChain_io_update_bits;
	wire clock_falling = ~clock;
	reg tdoReg;
	wire [3:0] currState = stateMachine_io_currState;
	wire _irChain_io_chainIn_update_T = currState == 4'hd;
	reg [4:0] activeInstruction;
	wire tapIsInTestLogicReset = currState == 4'hf;
	wire _io_dataChainOut_shift_T = currState == 4'h2;
	wire _GEN_2 = irChain_io_chainOut_data;
	JtagStateMachine stateMachine(
		.clock(stateMachine_clock),
		.reset(stateMachine_reset),
		.io_tms(stateMachine_io_tms),
		.io_currState(stateMachine_io_currState)
	);
	CaptureUpdateChain_2 irChain(
		.clock(irChain_clock),
		.reset(irChain_reset),
		.io_chainIn_shift(irChain_io_chainIn_shift),
		.io_chainIn_data(irChain_io_chainIn_data),
		.io_chainIn_capture(irChain_io_chainIn_capture),
		.io_chainIn_update(irChain_io_chainIn_update),
		.io_chainOut_data(irChain_io_chainOut_data),
		.io_update_bits(irChain_io_update_bits)
	);
	assign io_jtag_TDO_data = tdoReg;
	assign io_output_instruction = activeInstruction;
	assign io_output_tapIsInTestLogicReset = currState == 4'hf;
	assign io_dataChainOut_shift = currState == 4'h2;
	assign io_dataChainOut_data = io_jtag_TDI;
	assign io_dataChainOut_capture = currState == 4'h6;
	assign io_dataChainOut_update = currState == 4'h5;
	assign stateMachine_clock = clock;
	assign stateMachine_reset = io_control_jtag_reset;
	assign stateMachine_io_tms = io_jtag_TMS;
	assign irChain_clock = clock;
	assign irChain_reset = reset;
	assign irChain_io_chainIn_shift = currState == 4'ha;
	assign irChain_io_chainIn_data = io_jtag_TDI;
	assign irChain_io_chainIn_capture = currState == 4'he;
	assign irChain_io_chainIn_update = currState == 4'hd;
	always @(posedge clock_falling or posedge io_control_jtag_reset)
		if (io_control_jtag_reset)
			tdoReg <= 1'h0;
		else if (_io_dataChainOut_shift_T)
			tdoReg <= io_dataChainIn_data;
		else
			tdoReg <= _GEN_2;
	always @(posedge clock_falling or posedge io_control_jtag_reset)
		if (io_control_jtag_reset)
			activeInstruction <= 5'h01;
		else if (tapIsInTestLogicReset)
			activeInstruction <= 5'h01;
		else if (_irChain_io_chainIn_update_T)
			activeInstruction <= irChain_io_update_bits;
endmodule
module JtagBypassChain (
	clock,
	reset,
	io_chainIn_shift,
	io_chainIn_data,
	io_chainIn_capture,
	io_chainIn_update,
	io_chainOut_data
);
	input clock;
	input reset;
	input io_chainIn_shift;
	input io_chainIn_data;
	input io_chainIn_capture;
	input io_chainIn_update;
	output wire io_chainOut_data;
	reg reg_;
	wire _T_1 = ~(io_chainIn_capture & io_chainIn_update);
	wire _T_4 = _T_1 & ~(io_chainIn_capture & io_chainIn_shift);
	wire _T_7 = _T_4 & ~(io_chainIn_update & io_chainIn_shift);
	assign io_chainOut_data = reg_;
	always @(posedge clock)
		if (io_chainIn_capture)
			reg_ <= 1'h0;
		else if (io_chainIn_shift)
			reg_ <= io_chainIn_data;
endmodule
module DebugTransportModuleJTAG (
	io_jtag_clock,
	io_jtag_reset,
	io_dmi_req_ready,
	io_dmi_req_valid,
	io_dmi_req_bits_addr,
	io_dmi_req_bits_data,
	io_dmi_req_bits_op,
	io_dmi_resp_ready,
	io_dmi_resp_valid,
	io_dmi_resp_bits_data,
	io_dmi_resp_bits_resp,
	io_jtag_TMS,
	io_jtag_TDI,
	io_jtag_TDO_data
);
	input io_jtag_clock;
	input io_jtag_reset;
	input io_dmi_req_ready;
	output wire io_dmi_req_valid;
	output wire [6:0] io_dmi_req_bits_addr;
	output wire [31:0] io_dmi_req_bits_data;
	output wire [1:0] io_dmi_req_bits_op;
	output wire io_dmi_resp_ready;
	input io_dmi_resp_valid;
	input [31:0] io_dmi_resp_bits_data;
	input [1:0] io_dmi_resp_bits_resp;
	input io_jtag_TMS;
	input io_jtag_TDI;
	output wire io_jtag_TDO_data;
	wire dtmInfoChain_clock;
	wire dtmInfoChain_reset;
	wire dtmInfoChain_io_chainIn_shift;
	wire dtmInfoChain_io_chainIn_data;
	wire dtmInfoChain_io_chainIn_capture;
	wire dtmInfoChain_io_chainIn_update;
	wire dtmInfoChain_io_chainOut_data;
	wire [1:0] dtmInfoChain_io_capture_bits_dmiStatus;
	wire dtmInfoChain_io_update_valid;
	wire dtmInfoChain_io_update_bits_dmireset;
	wire dmiAccessChain_clock;
	wire dmiAccessChain_reset;
	wire dmiAccessChain_io_chainIn_shift;
	wire dmiAccessChain_io_chainIn_data;
	wire dmiAccessChain_io_chainIn_capture;
	wire dmiAccessChain_io_chainIn_update;
	wire dmiAccessChain_io_chainOut_data;
	wire [6:0] dmiAccessChain_io_capture_bits_addr;
	wire [31:0] dmiAccessChain_io_capture_bits_data;
	wire [1:0] dmiAccessChain_io_capture_bits_resp;
	wire dmiAccessChain_io_capture_capture;
	wire dmiAccessChain_io_update_valid;
	wire [6:0] dmiAccessChain_io_update_bits_addr;
	wire [31:0] dmiAccessChain_io_update_bits_data;
	wire [1:0] dmiAccessChain_io_update_bits_op;
	wire tapIO_idcodeChain_clock;
	wire tapIO_idcodeChain_reset;
	wire tapIO_idcodeChain_io_chainIn_shift;
	wire tapIO_idcodeChain_io_chainIn_data;
	wire tapIO_idcodeChain_io_chainIn_capture;
	wire tapIO_idcodeChain_io_chainIn_update;
	wire tapIO_idcodeChain_io_chainOut_data;
	wire tapIO_controllerInternal_clock;
	wire tapIO_controllerInternal_reset;
	wire tapIO_controllerInternal_io_jtag_TMS;
	wire tapIO_controllerInternal_io_jtag_TDI;
	wire tapIO_controllerInternal_io_jtag_TDO_data;
	wire tapIO_controllerInternal_io_control_jtag_reset;
	wire [4:0] tapIO_controllerInternal_io_output_instruction;
	wire tapIO_controllerInternal_io_output_tapIsInTestLogicReset;
	wire tapIO_controllerInternal_io_dataChainOut_shift;
	wire tapIO_controllerInternal_io_dataChainOut_data;
	wire tapIO_controllerInternal_io_dataChainOut_capture;
	wire tapIO_controllerInternal_io_dataChainOut_update;
	wire tapIO_controllerInternal_io_dataChainIn_data;
	wire tapIO_bypassChain_clock;
	wire tapIO_bypassChain_reset;
	wire tapIO_bypassChain_io_chainIn_shift;
	wire tapIO_bypassChain_io_chainIn_data;
	wire tapIO_bypassChain_io_chainIn_capture;
	wire tapIO_bypassChain_io_chainIn_update;
	wire tapIO_bypassChain_io_chainOut_data;
	reg busyReg;
	reg stickyBusyReg;
	reg stickyNonzeroRespReg;
	reg downgradeOpReg;
	reg [6:0] dmiReqReg_addr;
	reg [31:0] dmiReqReg_data;
	reg [1:0] dmiReqReg_op;
	reg dmiReqValidReg;
	wire _dmiStatus_T = stickyNonzeroRespReg | stickyBusyReg;
	wire _GEN_0 = io_dmi_req_valid | busyReg;
	wire _T_1 = io_dmi_resp_ready & io_dmi_resp_valid;
	wire busy = (busyReg & ~io_dmi_resp_valid) | stickyBusyReg;
	wire _downgradeOpReg_T = ~busy;
	wire nonzeroResp = stickyNonzeroRespReg | (io_dmi_resp_valid & (io_dmi_resp_bits_resp != 2'h0));
	wire _GEN_4 = (dmiAccessChain_io_capture_capture ? busy : stickyBusyReg);
	wire _GEN_5 = (dmiAccessChain_io_capture_capture ? nonzeroResp : stickyNonzeroRespReg);
	wire [6:0] _dmiAccessChain_io_capture_bits_T_addr = (io_dmi_resp_valid ? dmiReqReg_addr : 7'h00);
	wire [31:0] _dmiAccessChain_io_capture_bits_T_data = (io_dmi_resp_valid ? io_dmi_resp_bits_data : 32'h00000000);
	wire [1:0] _dmiAccessChain_io_capture_bits_T_resp = (io_dmi_resp_valid ? io_dmi_resp_bits_resp : 2'h0);
	wire _T_4 = io_dmi_req_ready & io_dmi_req_valid;
	wire _GEN_14 = (downgradeOpReg | (dmiAccessChain_io_update_bits_op == 2'h0) ? 1'h0 : 1'h1);
	wire _GEN_19 = (stickyBusyReg ? 1'h0 : _GEN_14);
	wire dmiReqValidCheck = dmiAccessChain_io_update_valid & _GEN_19;
	wire _T_8 = ~io_jtag_reset;
	wire _GEN_13 = (downgradeOpReg | (dmiAccessChain_io_update_bits_op == 2'h0) ? dmiReqValidReg : 1'h1);
	wire _io_dmi_resp_ready_T = dmiReqReg_op == 2'h2;
	wire _io_dmi_resp_ready_T_2 = dmiAccessChain_io_capture_capture & _downgradeOpReg_T;
	wire [31:0] _GEN_1 = 32'h00000001 % 32'h00000002;
	wire [1:0] _tapIO_T = _GEN_1[1:0];
	wire tapIO_icodeSelects_0 = tapIO_controllerInternal_io_output_instruction == 5'h01;
	wire tapIO_icodeSelects_0_1 = tapIO_controllerInternal_io_output_instruction == 5'h10;
	wire tapIO_icodeSelects_0_2 = tapIO_controllerInternal_io_output_instruction == 5'h11;
	wire _GEN_28 = (tapIO_icodeSelects_0_2 ? dmiAccessChain_io_chainOut_data : tapIO_bypassChain_io_chainOut_data);
	wire _GEN_32 = (tapIO_icodeSelects_0_1 ? dtmInfoChain_io_chainOut_data : _GEN_28);
	wire tapIO_output_tapIsInTestLogicReset = tapIO_controllerInternal_io_output_tapIsInTestLogicReset;
	CaptureUpdateChain dtmInfoChain(
		.clock(dtmInfoChain_clock),
		.reset(dtmInfoChain_reset),
		.io_chainIn_shift(dtmInfoChain_io_chainIn_shift),
		.io_chainIn_data(dtmInfoChain_io_chainIn_data),
		.io_chainIn_capture(dtmInfoChain_io_chainIn_capture),
		.io_chainIn_update(dtmInfoChain_io_chainIn_update),
		.io_chainOut_data(dtmInfoChain_io_chainOut_data),
		.io_capture_bits_dmiStatus(dtmInfoChain_io_capture_bits_dmiStatus),
		.io_update_valid(dtmInfoChain_io_update_valid),
		.io_update_bits_dmireset(dtmInfoChain_io_update_bits_dmireset)
	);
	CaptureUpdateChain_1 dmiAccessChain(
		.clock(dmiAccessChain_clock),
		.reset(dmiAccessChain_reset),
		.io_chainIn_shift(dmiAccessChain_io_chainIn_shift),
		.io_chainIn_data(dmiAccessChain_io_chainIn_data),
		.io_chainIn_capture(dmiAccessChain_io_chainIn_capture),
		.io_chainIn_update(dmiAccessChain_io_chainIn_update),
		.io_chainOut_data(dmiAccessChain_io_chainOut_data),
		.io_capture_bits_addr(dmiAccessChain_io_capture_bits_addr),
		.io_capture_bits_data(dmiAccessChain_io_capture_bits_data),
		.io_capture_bits_resp(dmiAccessChain_io_capture_bits_resp),
		.io_capture_capture(dmiAccessChain_io_capture_capture),
		.io_update_valid(dmiAccessChain_io_update_valid),
		.io_update_bits_addr(dmiAccessChain_io_update_bits_addr),
		.io_update_bits_data(dmiAccessChain_io_update_bits_data),
		.io_update_bits_op(dmiAccessChain_io_update_bits_op)
	);
	CaptureChain tapIO_idcodeChain(
		.clock(tapIO_idcodeChain_clock),
		.reset(tapIO_idcodeChain_reset),
		.io_chainIn_shift(tapIO_idcodeChain_io_chainIn_shift),
		.io_chainIn_data(tapIO_idcodeChain_io_chainIn_data),
		.io_chainIn_capture(tapIO_idcodeChain_io_chainIn_capture),
		.io_chainIn_update(tapIO_idcodeChain_io_chainIn_update),
		.io_chainOut_data(tapIO_idcodeChain_io_chainOut_data)
	);
	JtagTapController tapIO_controllerInternal(
		.clock(tapIO_controllerInternal_clock),
		.reset(tapIO_controllerInternal_reset),
		.io_jtag_TMS(tapIO_controllerInternal_io_jtag_TMS),
		.io_jtag_TDI(tapIO_controllerInternal_io_jtag_TDI),
		.io_jtag_TDO_data(tapIO_controllerInternal_io_jtag_TDO_data),
		.io_control_jtag_reset(tapIO_controllerInternal_io_control_jtag_reset),
		.io_output_instruction(tapIO_controllerInternal_io_output_instruction),
		.io_output_tapIsInTestLogicReset(tapIO_controllerInternal_io_output_tapIsInTestLogicReset),
		.io_dataChainOut_shift(tapIO_controllerInternal_io_dataChainOut_shift),
		.io_dataChainOut_data(tapIO_controllerInternal_io_dataChainOut_data),
		.io_dataChainOut_capture(tapIO_controllerInternal_io_dataChainOut_capture),
		.io_dataChainOut_update(tapIO_controllerInternal_io_dataChainOut_update),
		.io_dataChainIn_data(tapIO_controllerInternal_io_dataChainIn_data)
	);
	JtagBypassChain tapIO_bypassChain(
		.clock(tapIO_bypassChain_clock),
		.reset(tapIO_bypassChain_reset),
		.io_chainIn_shift(tapIO_bypassChain_io_chainIn_shift),
		.io_chainIn_data(tapIO_bypassChain_io_chainIn_data),
		.io_chainIn_capture(tapIO_bypassChain_io_chainIn_capture),
		.io_chainIn_update(tapIO_bypassChain_io_chainIn_update),
		.io_chainOut_data(tapIO_bypassChain_io_chainOut_data)
	);
	assign io_dmi_req_valid = dmiReqValidReg;
	assign io_dmi_req_bits_addr = dmiReqReg_addr;
	assign io_dmi_req_bits_data = dmiReqReg_data;
	assign io_dmi_req_bits_op = dmiReqReg_op;
	assign io_dmi_resp_ready = (_io_dmi_resp_ready_T ? io_dmi_resp_valid : _io_dmi_resp_ready_T_2);
	assign io_jtag_TDO_data = tapIO_controllerInternal_io_jtag_TDO_data;
	assign dtmInfoChain_clock = io_jtag_clock;
	assign dtmInfoChain_reset = io_jtag_reset;
	assign dtmInfoChain_io_chainIn_shift = tapIO_icodeSelects_0_1 & tapIO_controllerInternal_io_dataChainOut_shift;
	assign dtmInfoChain_io_chainIn_data = tapIO_icodeSelects_0_1 & tapIO_controllerInternal_io_dataChainOut_data;
	assign dtmInfoChain_io_chainIn_capture = tapIO_icodeSelects_0_1 & tapIO_controllerInternal_io_dataChainOut_capture;
	assign dtmInfoChain_io_chainIn_update = tapIO_icodeSelects_0_1 & tapIO_controllerInternal_io_dataChainOut_update;
	assign dtmInfoChain_io_capture_bits_dmiStatus = {stickyNonzeroRespReg, _dmiStatus_T};
	assign dmiAccessChain_clock = io_jtag_clock;
	assign dmiAccessChain_reset = io_jtag_reset;
	assign dmiAccessChain_io_chainIn_shift = tapIO_icodeSelects_0_2 & tapIO_controllerInternal_io_dataChainOut_shift;
	assign dmiAccessChain_io_chainIn_data = tapIO_icodeSelects_0_2 & tapIO_controllerInternal_io_dataChainOut_data;
	assign dmiAccessChain_io_chainIn_capture = tapIO_icodeSelects_0_2 & tapIO_controllerInternal_io_dataChainOut_capture;
	assign dmiAccessChain_io_chainIn_update = tapIO_icodeSelects_0_2 & tapIO_controllerInternal_io_dataChainOut_update;
	assign dmiAccessChain_io_capture_bits_addr = (busy ? 7'h00 : _dmiAccessChain_io_capture_bits_T_addr);
	assign dmiAccessChain_io_capture_bits_data = (busy ? 32'h00000000 : _dmiAccessChain_io_capture_bits_T_data);
	assign dmiAccessChain_io_capture_bits_resp = (busy ? 2'h3 : _dmiAccessChain_io_capture_bits_T_resp);
	assign tapIO_idcodeChain_clock = io_jtag_clock;
	assign tapIO_idcodeChain_reset = io_jtag_reset;
	assign tapIO_idcodeChain_io_chainIn_shift = tapIO_icodeSelects_0 & tapIO_controllerInternal_io_dataChainOut_shift;
	assign tapIO_idcodeChain_io_chainIn_data = tapIO_icodeSelects_0 & tapIO_controllerInternal_io_dataChainOut_data;
	assign tapIO_idcodeChain_io_chainIn_capture = tapIO_icodeSelects_0 & tapIO_controllerInternal_io_dataChainOut_capture;
	assign tapIO_idcodeChain_io_chainIn_update = tapIO_icodeSelects_0 & tapIO_controllerInternal_io_dataChainOut_update;
	assign tapIO_controllerInternal_clock = io_jtag_clock;
	assign tapIO_controllerInternal_reset = io_jtag_reset;
	assign tapIO_controllerInternal_io_jtag_TMS = io_jtag_TMS;
	assign tapIO_controllerInternal_io_jtag_TDI = io_jtag_TDI;
	assign tapIO_controllerInternal_io_control_jtag_reset = io_jtag_reset;
	assign tapIO_controllerInternal_io_dataChainIn_data = (tapIO_icodeSelects_0 ? tapIO_idcodeChain_io_chainOut_data : _GEN_32);
	assign tapIO_bypassChain_clock = io_jtag_clock;
	assign tapIO_bypassChain_reset = io_jtag_reset;
	assign tapIO_bypassChain_io_chainIn_shift = tapIO_controllerInternal_io_dataChainOut_shift;
	assign tapIO_bypassChain_io_chainIn_data = tapIO_controllerInternal_io_dataChainOut_data;
	assign tapIO_bypassChain_io_chainIn_capture = tapIO_controllerInternal_io_dataChainOut_capture;
	assign tapIO_bypassChain_io_chainIn_update = tapIO_controllerInternal_io_dataChainOut_update;
	always @(posedge io_jtag_clock) begin
		if (dmiAccessChain_io_update_valid)
			if (!stickyBusyReg)
				if (downgradeOpReg | (dmiAccessChain_io_update_bits_op == 2'h0))
					dmiReqReg_addr <= 7'h00;
				else
					dmiReqReg_addr <= dmiAccessChain_io_update_bits_addr;
		if (dmiAccessChain_io_update_valid)
			if (!stickyBusyReg)
				if (downgradeOpReg | (dmiAccessChain_io_update_bits_op == 2'h0))
					dmiReqReg_data <= 32'h00000000;
				else
					dmiReqReg_data <= dmiAccessChain_io_update_bits_data;
		if (dmiAccessChain_io_update_valid)
			if (!stickyBusyReg)
				if (downgradeOpReg | (dmiAccessChain_io_update_bits_op == 2'h0))
					dmiReqReg_op <= 2'h0;
				else
					dmiReqReg_op <= dmiAccessChain_io_update_bits_op;
	end
	always @(posedge io_jtag_clock or posedge io_jtag_reset)
		if (io_jtag_reset)
			busyReg <= 1'h0;
		else if (tapIO_output_tapIsInTestLogicReset)
			busyReg <= 1'h0;
		else if (_T_1)
			busyReg <= 1'h0;
		else
			busyReg <= _GEN_0;
	always @(posedge io_jtag_clock or posedge io_jtag_reset)
		if (io_jtag_reset)
			stickyBusyReg <= 1'h0;
		else if (tapIO_output_tapIsInTestLogicReset)
			stickyBusyReg <= 1'h0;
		else if (dtmInfoChain_io_update_valid) begin
			if (dtmInfoChain_io_update_bits_dmireset)
				stickyBusyReg <= 1'h0;
			else
				stickyBusyReg <= _GEN_4;
		end
		else
			stickyBusyReg <= _GEN_4;
	always @(posedge io_jtag_clock or posedge io_jtag_reset)
		if (io_jtag_reset)
			stickyNonzeroRespReg <= 1'h0;
		else if (tapIO_output_tapIsInTestLogicReset)
			stickyNonzeroRespReg <= 1'h0;
		else if (dtmInfoChain_io_update_valid) begin
			if (dtmInfoChain_io_update_bits_dmireset)
				stickyNonzeroRespReg <= 1'h0;
			else
				stickyNonzeroRespReg <= _GEN_5;
		end
		else
			stickyNonzeroRespReg <= _GEN_5;
	always @(posedge io_jtag_clock or posedge io_jtag_reset)
		if (io_jtag_reset)
			downgradeOpReg <= 1'h0;
		else if (tapIO_output_tapIsInTestLogicReset)
			downgradeOpReg <= 1'h0;
		else if (dmiAccessChain_io_capture_capture)
			downgradeOpReg <= ~busy & nonzeroResp;
		else if (dmiAccessChain_io_update_valid)
			downgradeOpReg <= 1'h0;
	always @(posedge io_jtag_clock or posedge io_jtag_reset)
		if (io_jtag_reset)
			dmiReqValidReg <= 1'h0;
		else if (tapIO_output_tapIsInTestLogicReset)
			dmiReqValidReg <= 1'h0;
		else if (_T_4)
			dmiReqValidReg <= 1'h0;
		else if (dmiAccessChain_io_update_valid)
			if (!stickyBusyReg)
				dmiReqValidReg <= _GEN_13;
endmodule
module DigitalTop (
	clock,
	reset,
	auto_implicitClockGrouper_out_clock,
	auto_implicitClockGrouper_out_reset,
	auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock,
	auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset,
	auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock,
	auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset,
	auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock,
	auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset,
	auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock,
	auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset,
	auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock,
	auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset,
	auto_subsystem_cbus_fixedClockNode_out_clock,
	auto_subsystem_cbus_fixedClockNode_out_reset,
	custom_boot,
	serial_tl_clock,
	serial_tl_bits_in_ready,
	serial_tl_bits_in_valid,
	serial_tl_bits_in_bits,
	serial_tl_bits_out_ready,
	serial_tl_bits_out_valid,
	serial_tl_bits_out_bits,
	resetctrl_hartIsInReset_0,
	debug_clock,
	debug_reset,
	debug_systemjtag_jtag_TCK,
	debug_systemjtag_jtag_TMS,
	debug_systemjtag_jtag_TDI,
	debug_systemjtag_jtag_TDO_data,
	debug_systemjtag_reset,
	debug_dmactive,
	debug_dmactiveAck,
	uart_0_txd,
	uart_0_rxd
);
	input clock;
	input reset;
	output wire auto_implicitClockGrouper_out_clock;
	output wire auto_implicitClockGrouper_out_reset;
	input auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock;
	input auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset;
	input auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock;
	input auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset;
	input auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock;
	input auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset;
	input auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock;
	input auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset;
	input auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock;
	input auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset;
	output wire auto_subsystem_cbus_fixedClockNode_out_clock;
	output wire auto_subsystem_cbus_fixedClockNode_out_reset;
	input custom_boot;
	output wire serial_tl_clock;
	output wire serial_tl_bits_in_ready;
	input serial_tl_bits_in_valid;
	input [31:0] serial_tl_bits_in_bits;
	input serial_tl_bits_out_ready;
	output wire serial_tl_bits_out_valid;
	output wire [31:0] serial_tl_bits_out_bits;
	input resetctrl_hartIsInReset_0;
	input debug_clock;
	input debug_reset;
	input debug_systemjtag_jtag_TCK;
	input debug_systemjtag_jtag_TMS;
	input debug_systemjtag_jtag_TDI;
	output wire debug_systemjtag_jtag_TDO_data;
	input debug_systemjtag_reset;
	output wire debug_dmactive;
	input debug_dmactiveAck;
	output wire uart_0_txd;
	input uart_0_rxd;
	wire ibus_auto_int_bus_int_in_0;
	wire ibus_auto_int_bus_int_out_0;
	wire subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_ready;
	wire subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_valid;
	wire [2:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode;
	wire [2:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param;
	wire [3:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size;
	wire subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source;
	wire [31:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address;
	wire [3:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask;
	wire [31:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data;
	wire subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_corrupt;
	wire subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_ready;
	wire subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_valid;
	wire [2:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode;
	wire [1:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param;
	wire [3:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size;
	wire subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source;
	wire subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink;
	wire subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied;
	wire [31:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data;
	wire subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt;
	wire subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready;
	wire subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid;
	wire [2:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode;
	wire [2:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param;
	wire [3:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size;
	wire subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source;
	wire [31:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address;
	wire [3:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask;
	wire [31:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data;
	wire subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_corrupt;
	wire subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready;
	wire subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid;
	wire [2:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode;
	wire [1:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param;
	wire [3:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size;
	wire subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink;
	wire subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied;
	wire [31:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data;
	wire subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt;
	wire subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready;
	wire subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid;
	wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode;
	wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param;
	wire [3:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size;
	wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source;
	wire [31:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address;
	wire [3:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask;
	wire [31:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data;
	wire subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt;
	wire subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready;
	wire subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid;
	wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode;
	wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param;
	wire [3:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size;
	wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source;
	wire subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink;
	wire subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied;
	wire [31:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data;
	wire subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt;
	wire subsystem_sbus_auto_fixedClockNode_out_1_clock;
	wire subsystem_sbus_auto_fixedClockNode_out_1_reset;
	wire subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock;
	wire subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset;
	wire subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_ready;
	wire subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_valid;
	wire [2:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode;
	wire [2:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_param;
	wire [1:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size;
	wire [7:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source;
	wire [30:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address;
	wire [3:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask;
	wire [31:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data;
	wire subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_corrupt;
	wire subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_ready;
	wire subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_valid;
	wire [2:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode;
	wire [1:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size;
	wire [7:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source;
	wire [31:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data;
	wire subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_ready;
	wire subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_valid;
	wire [2:0] subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_opcode;
	wire [2:0] subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_param;
	wire [2:0] subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_size;
	wire [2:0] subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_source;
	wire [28:0] subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_address;
	wire [7:0] subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_mask;
	wire [63:0] subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_data;
	wire subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_corrupt;
	wire subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_ready;
	wire subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_valid;
	wire [2:0] subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_opcode;
	wire [1:0] subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_param;
	wire [2:0] subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_size;
	wire [2:0] subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_source;
	wire subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_sink;
	wire subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_denied;
	wire [63:0] subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_data;
	wire subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_corrupt;
	wire subsystem_pbus_auto_fixedClockNode_out_clock;
	wire subsystem_pbus_auto_fixedClockNode_out_reset;
	wire subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock;
	wire subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset;
	wire subsystem_pbus_auto_bus_xing_in_a_ready;
	wire subsystem_pbus_auto_bus_xing_in_a_valid;
	wire [2:0] subsystem_pbus_auto_bus_xing_in_a_bits_opcode;
	wire [2:0] subsystem_pbus_auto_bus_xing_in_a_bits_param;
	wire [2:0] subsystem_pbus_auto_bus_xing_in_a_bits_size;
	wire [2:0] subsystem_pbus_auto_bus_xing_in_a_bits_source;
	wire [30:0] subsystem_pbus_auto_bus_xing_in_a_bits_address;
	wire [3:0] subsystem_pbus_auto_bus_xing_in_a_bits_mask;
	wire [31:0] subsystem_pbus_auto_bus_xing_in_a_bits_data;
	wire subsystem_pbus_auto_bus_xing_in_a_bits_corrupt;
	wire subsystem_pbus_auto_bus_xing_in_d_ready;
	wire subsystem_pbus_auto_bus_xing_in_d_valid;
	wire [2:0] subsystem_pbus_auto_bus_xing_in_d_bits_opcode;
	wire [1:0] subsystem_pbus_auto_bus_xing_in_d_bits_param;
	wire [2:0] subsystem_pbus_auto_bus_xing_in_d_bits_size;
	wire [2:0] subsystem_pbus_auto_bus_xing_in_d_bits_source;
	wire subsystem_pbus_auto_bus_xing_in_d_bits_sink;
	wire subsystem_pbus_auto_bus_xing_in_d_bits_denied;
	wire [31:0] subsystem_pbus_auto_bus_xing_in_d_bits_data;
	wire subsystem_pbus_auto_bus_xing_in_d_bits_corrupt;
	wire subsystem_pbus_clock;
	wire subsystem_pbus_reset;
	wire subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_ready;
	wire subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_valid;
	wire [2:0] subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_opcode;
	wire [2:0] subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_param;
	wire [3:0] subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_size;
	wire subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_source;
	wire [31:0] subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_address;
	wire [3:0] subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_mask;
	wire [31:0] subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_data;
	wire subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_corrupt;
	wire subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_ready;
	wire subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_valid;
	wire [2:0] subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_opcode;
	wire [1:0] subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_param;
	wire [3:0] subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_size;
	wire subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_source;
	wire subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_sink;
	wire subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_denied;
	wire [31:0] subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_data;
	wire subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_corrupt;
	wire subsystem_fbus_auto_fixedClockNode_out_clock;
	wire subsystem_fbus_auto_fixedClockNode_out_reset;
	wire subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock;
	wire subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset;
	wire subsystem_fbus_auto_bus_xing_out_a_ready;
	wire subsystem_fbus_auto_bus_xing_out_a_valid;
	wire [2:0] subsystem_fbus_auto_bus_xing_out_a_bits_opcode;
	wire [2:0] subsystem_fbus_auto_bus_xing_out_a_bits_param;
	wire [3:0] subsystem_fbus_auto_bus_xing_out_a_bits_size;
	wire subsystem_fbus_auto_bus_xing_out_a_bits_source;
	wire [31:0] subsystem_fbus_auto_bus_xing_out_a_bits_address;
	wire [3:0] subsystem_fbus_auto_bus_xing_out_a_bits_mask;
	wire [31:0] subsystem_fbus_auto_bus_xing_out_a_bits_data;
	wire subsystem_fbus_auto_bus_xing_out_a_bits_corrupt;
	wire subsystem_fbus_auto_bus_xing_out_d_ready;
	wire subsystem_fbus_auto_bus_xing_out_d_valid;
	wire [2:0] subsystem_fbus_auto_bus_xing_out_d_bits_opcode;
	wire [1:0] subsystem_fbus_auto_bus_xing_out_d_bits_param;
	wire [3:0] subsystem_fbus_auto_bus_xing_out_d_bits_size;
	wire subsystem_fbus_auto_bus_xing_out_d_bits_sink;
	wire subsystem_fbus_auto_bus_xing_out_d_bits_denied;
	wire [31:0] subsystem_fbus_auto_bus_xing_out_d_bits_data;
	wire subsystem_fbus_auto_bus_xing_out_d_bits_corrupt;
	wire subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_ready;
	wire subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_opcode;
	wire [2:0] subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_param;
	wire [1:0] subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_size;
	wire [7:0] subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_source;
	wire [20:0] subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_address;
	wire [3:0] subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_mask;
	wire [31:0] subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_data;
	wire subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_corrupt;
	wire subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_ready;
	wire subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_opcode;
	wire [1:0] subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_size;
	wire [7:0] subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_source;
	wire [31:0] subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_data;
	wire subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_ready;
	wire subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_opcode;
	wire [2:0] subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_param;
	wire [1:0] subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_size;
	wire [7:0] subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_source;
	wire [20:0] subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_address;
	wire [3:0] subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_mask;
	wire [31:0] subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_data;
	wire subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_corrupt;
	wire subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_ready;
	wire subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_opcode;
	wire [1:0] subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_size;
	wire [7:0] subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_source;
	wire [31:0] subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_data;
	wire subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_ready;
	wire subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode;
	wire [2:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_param;
	wire [1:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_size;
	wire [7:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_source;
	wire [16:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_address;
	wire [3:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_mask;
	wire subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt;
	wire subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_ready;
	wire subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_valid;
	wire [1:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_size;
	wire [7:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_source;
	wire [31:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_data;
	wire subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_ready;
	wire subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_opcode;
	wire [2:0] subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_param;
	wire [2:0] subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_size;
	wire [2:0] subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_source;
	wire [31:0] subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_address;
	wire [3:0] subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_mask;
	wire [31:0] subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_data;
	wire subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_ready;
	wire subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_opcode;
	wire [1:0] subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_param;
	wire [2:0] subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_size;
	wire [2:0] subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_source;
	wire subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_sink;
	wire subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_denied;
	wire [31:0] subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_data;
	wire subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_corrupt;
	wire subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_ready;
	wire subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_opcode;
	wire [2:0] subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_param;
	wire [1:0] subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_size;
	wire [7:0] subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_source;
	wire [11:0] subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_address;
	wire [3:0] subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_mask;
	wire [31:0] subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_data;
	wire subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_corrupt;
	wire subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_ready;
	wire subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_bits_opcode;
	wire [1:0] subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_bits_size;
	wire [7:0] subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_bits_source;
	wire [31:0] subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_bits_data;
	wire subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_ready;
	wire subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_opcode;
	wire [2:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_param;
	wire [1:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_size;
	wire [7:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_source;
	wire [25:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_address;
	wire [3:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_mask;
	wire [31:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_data;
	wire subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_corrupt;
	wire subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_ready;
	wire subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_opcode;
	wire [1:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_size;
	wire [7:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_source;
	wire [31:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_data;
	wire subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_ready;
	wire subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_opcode;
	wire [2:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_param;
	wire [1:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_size;
	wire [7:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_source;
	wire [27:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_address;
	wire [3:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_mask;
	wire [31:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_data;
	wire subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_corrupt;
	wire subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_ready;
	wire subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_opcode;
	wire [1:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_size;
	wire [7:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_source;
	wire [31:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_data;
	wire subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready;
	wire subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode;
	wire [2:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param;
	wire [2:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size;
	wire [2:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source;
	wire [30:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address;
	wire [3:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask;
	wire [31:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data;
	wire subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_corrupt;
	wire subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready;
	wire subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid;
	wire [2:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode;
	wire [1:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_param;
	wire [2:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size;
	wire [2:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source;
	wire subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_sink;
	wire subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied;
	wire [31:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data;
	wire subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt;
	wire subsystem_cbus_auto_fixedClockNode_out_4_clock;
	wire subsystem_cbus_auto_fixedClockNode_out_4_reset;
	wire subsystem_cbus_auto_fixedClockNode_out_3_clock;
	wire subsystem_cbus_auto_fixedClockNode_out_3_reset;
	wire subsystem_cbus_auto_fixedClockNode_out_2_clock;
	wire subsystem_cbus_auto_fixedClockNode_out_2_reset;
	wire subsystem_cbus_auto_fixedClockNode_out_0_clock;
	wire subsystem_cbus_auto_fixedClockNode_out_0_reset;
	wire subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock;
	wire subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset;
	wire subsystem_cbus_auto_bus_xing_in_a_ready;
	wire subsystem_cbus_auto_bus_xing_in_a_valid;
	wire [2:0] subsystem_cbus_auto_bus_xing_in_a_bits_opcode;
	wire [2:0] subsystem_cbus_auto_bus_xing_in_a_bits_param;
	wire [3:0] subsystem_cbus_auto_bus_xing_in_a_bits_size;
	wire [1:0] subsystem_cbus_auto_bus_xing_in_a_bits_source;
	wire [31:0] subsystem_cbus_auto_bus_xing_in_a_bits_address;
	wire [3:0] subsystem_cbus_auto_bus_xing_in_a_bits_mask;
	wire [31:0] subsystem_cbus_auto_bus_xing_in_a_bits_data;
	wire subsystem_cbus_auto_bus_xing_in_a_bits_corrupt;
	wire subsystem_cbus_auto_bus_xing_in_d_ready;
	wire subsystem_cbus_auto_bus_xing_in_d_valid;
	wire [2:0] subsystem_cbus_auto_bus_xing_in_d_bits_opcode;
	wire [1:0] subsystem_cbus_auto_bus_xing_in_d_bits_param;
	wire [3:0] subsystem_cbus_auto_bus_xing_in_d_bits_size;
	wire [1:0] subsystem_cbus_auto_bus_xing_in_d_bits_source;
	wire subsystem_cbus_auto_bus_xing_in_d_bits_sink;
	wire subsystem_cbus_auto_bus_xing_in_d_bits_denied;
	wire [31:0] subsystem_cbus_auto_bus_xing_in_d_bits_data;
	wire subsystem_cbus_auto_bus_xing_in_d_bits_corrupt;
	wire subsystem_cbus_custom_boot;
	wire subsystem_cbus_clock;
	wire subsystem_cbus_reset;
	wire tile_prci_domain_auto_intsink_in_sync_0;
	wire tile_prci_domain_auto_tile_reset_domain_tile_hartid_in;
	wire tile_prci_domain_auto_int_out_clock_xing_out_2_sync_0;
	wire tile_prci_domain_auto_int_out_clock_xing_out_1_sync_0;
	wire tile_prci_domain_auto_int_out_clock_xing_out_0_sync_0;
	wire tile_prci_domain_auto_int_in_clock_xing_in_1_sync_0;
	wire tile_prci_domain_auto_int_in_clock_xing_in_0_sync_0;
	wire tile_prci_domain_auto_int_in_clock_xing_in_0_sync_1;
	wire tile_prci_domain_auto_tl_slave_clock_xing_in_a_ready;
	wire tile_prci_domain_auto_tl_slave_clock_xing_in_a_valid;
	wire [2:0] tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_opcode;
	wire [2:0] tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_param;
	wire [2:0] tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_size;
	wire [2:0] tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_source;
	wire [31:0] tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_address;
	wire [3:0] tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_mask;
	wire [31:0] tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_data;
	wire tile_prci_domain_auto_tl_slave_clock_xing_in_d_ready;
	wire tile_prci_domain_auto_tl_slave_clock_xing_in_d_valid;
	wire [2:0] tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_opcode;
	wire [1:0] tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_param;
	wire [2:0] tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_size;
	wire [2:0] tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_source;
	wire tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_sink;
	wire tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_denied;
	wire [31:0] tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_data;
	wire tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_corrupt;
	wire tile_prci_domain_auto_tl_master_clock_xing_out_a_ready;
	wire tile_prci_domain_auto_tl_master_clock_xing_out_a_valid;
	wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_opcode;
	wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_param;
	wire [3:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_size;
	wire tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_source;
	wire [31:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_address;
	wire [3:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_mask;
	wire [31:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_data;
	wire tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_corrupt;
	wire tile_prci_domain_auto_tl_master_clock_xing_out_d_ready;
	wire tile_prci_domain_auto_tl_master_clock_xing_out_d_valid;
	wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_opcode;
	wire [1:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_param;
	wire [3:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_size;
	wire tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_source;
	wire tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_sink;
	wire tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_denied;
	wire [31:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_data;
	wire tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_corrupt;
	wire tile_prci_domain_auto_tap_clock_in_clock;
	wire tile_prci_domain_auto_tap_clock_in_reset;
	wire plicDomainWrapper_auto_plic_int_in_0;
	wire plicDomainWrapper_auto_plic_int_out_0;
	wire plicDomainWrapper_auto_plic_in_a_ready;
	wire plicDomainWrapper_auto_plic_in_a_valid;
	wire [2:0] plicDomainWrapper_auto_plic_in_a_bits_opcode;
	wire [2:0] plicDomainWrapper_auto_plic_in_a_bits_param;
	wire [1:0] plicDomainWrapper_auto_plic_in_a_bits_size;
	wire [7:0] plicDomainWrapper_auto_plic_in_a_bits_source;
	wire [27:0] plicDomainWrapper_auto_plic_in_a_bits_address;
	wire [3:0] plicDomainWrapper_auto_plic_in_a_bits_mask;
	wire [31:0] plicDomainWrapper_auto_plic_in_a_bits_data;
	wire plicDomainWrapper_auto_plic_in_a_bits_corrupt;
	wire plicDomainWrapper_auto_plic_in_d_ready;
	wire plicDomainWrapper_auto_plic_in_d_valid;
	wire [2:0] plicDomainWrapper_auto_plic_in_d_bits_opcode;
	wire [1:0] plicDomainWrapper_auto_plic_in_d_bits_size;
	wire [7:0] plicDomainWrapper_auto_plic_in_d_bits_source;
	wire [31:0] plicDomainWrapper_auto_plic_in_d_bits_data;
	wire plicDomainWrapper_auto_clock_in_clock;
	wire plicDomainWrapper_auto_clock_in_reset;
	wire clint_clock;
	wire clint_reset;
	wire clint_auto_int_out_0;
	wire clint_auto_int_out_1;
	wire clint_auto_in_a_ready;
	wire clint_auto_in_a_valid;
	wire [2:0] clint_auto_in_a_bits_opcode;
	wire [2:0] clint_auto_in_a_bits_param;
	wire [1:0] clint_auto_in_a_bits_size;
	wire [7:0] clint_auto_in_a_bits_source;
	wire [25:0] clint_auto_in_a_bits_address;
	wire [3:0] clint_auto_in_a_bits_mask;
	wire [31:0] clint_auto_in_a_bits_data;
	wire clint_auto_in_a_bits_corrupt;
	wire clint_auto_in_d_ready;
	wire clint_auto_in_d_valid;
	wire [2:0] clint_auto_in_d_bits_opcode;
	wire [1:0] clint_auto_in_d_bits_size;
	wire [7:0] clint_auto_in_d_bits_source;
	wire [31:0] clint_auto_in_d_bits_data;
	wire clint_io_rtcTick;
	wire debug_1_auto_dmInner_dmInner_tl_in_a_ready;
	wire debug_1_auto_dmInner_dmInner_tl_in_a_valid;
	wire [2:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_opcode;
	wire [2:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_param;
	wire [1:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_size;
	wire [7:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_source;
	wire [11:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_address;
	wire [3:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_mask;
	wire [31:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_data;
	wire debug_1_auto_dmInner_dmInner_tl_in_a_bits_corrupt;
	wire debug_1_auto_dmInner_dmInner_tl_in_d_ready;
	wire debug_1_auto_dmInner_dmInner_tl_in_d_valid;
	wire [2:0] debug_1_auto_dmInner_dmInner_tl_in_d_bits_opcode;
	wire [1:0] debug_1_auto_dmInner_dmInner_tl_in_d_bits_size;
	wire [7:0] debug_1_auto_dmInner_dmInner_tl_in_d_bits_source;
	wire [31:0] debug_1_auto_dmInner_dmInner_tl_in_d_bits_data;
	wire debug_1_auto_dmOuter_intsource_out_sync_0;
	wire debug_1_io_debug_clock;
	wire debug_1_io_debug_reset;
	wire debug_1_io_ctrl_dmactive;
	wire debug_1_io_ctrl_dmactiveAck;
	wire debug_1_io_dmi_dmi_req_ready;
	wire debug_1_io_dmi_dmi_req_valid;
	wire [6:0] debug_1_io_dmi_dmi_req_bits_addr;
	wire [31:0] debug_1_io_dmi_dmi_req_bits_data;
	wire [1:0] debug_1_io_dmi_dmi_req_bits_op;
	wire debug_1_io_dmi_dmi_resp_ready;
	wire debug_1_io_dmi_dmi_resp_valid;
	wire [31:0] debug_1_io_dmi_dmi_resp_bits_data;
	wire [1:0] debug_1_io_dmi_dmi_resp_bits_resp;
	wire debug_1_io_dmi_dmiClock;
	wire debug_1_io_dmi_dmiReset;
	wire debug_1_io_hartIsInReset_0;
	wire xbar_auto_int_in_0;
	wire xbar_auto_int_out_0;
	wire xbar_1_auto_int_in_0;
	wire xbar_1_auto_int_out_0;
	wire xbar_2_auto_int_in_0;
	wire xbar_2_auto_int_out_0;
	wire tileHartIdNexusNode_auto_out;
	wire intsource_clock;
	wire intsource_reset;
	wire intsource_auto_in_0;
	wire intsource_auto_in_1;
	wire intsource_auto_out_sync_0;
	wire intsource_auto_out_sync_1;
	wire intsource_1_clock;
	wire intsource_1_reset;
	wire intsource_1_auto_in_0;
	wire intsource_1_auto_out_sync_0;
	wire intsink_1_auto_in_sync_0;
	wire intsink_1_auto_out_0;
	wire intsink_2_auto_in_sync_0;
	wire intsink_2_auto_out_0;
	wire intsink_3_auto_in_sync_0;
	wire intsink_3_auto_out_0;
	wire bootROMDomainWrapper_auto_bootrom_in_a_ready;
	wire bootROMDomainWrapper_auto_bootrom_in_a_valid;
	wire [2:0] bootROMDomainWrapper_auto_bootrom_in_a_bits_opcode;
	wire [2:0] bootROMDomainWrapper_auto_bootrom_in_a_bits_param;
	wire [1:0] bootROMDomainWrapper_auto_bootrom_in_a_bits_size;
	wire [7:0] bootROMDomainWrapper_auto_bootrom_in_a_bits_source;
	wire [16:0] bootROMDomainWrapper_auto_bootrom_in_a_bits_address;
	wire [3:0] bootROMDomainWrapper_auto_bootrom_in_a_bits_mask;
	wire bootROMDomainWrapper_auto_bootrom_in_a_bits_corrupt;
	wire bootROMDomainWrapper_auto_bootrom_in_d_ready;
	wire bootROMDomainWrapper_auto_bootrom_in_d_valid;
	wire [1:0] bootROMDomainWrapper_auto_bootrom_in_d_bits_size;
	wire [7:0] bootROMDomainWrapper_auto_bootrom_in_d_bits_source;
	wire [31:0] bootROMDomainWrapper_auto_bootrom_in_d_bits_data;
	wire bootROMDomainWrapper_auto_clock_in_clock;
	wire bootROMDomainWrapper_auto_clock_in_reset;
	wire domain_auto_serdesser_client_out_a_ready;
	wire domain_auto_serdesser_client_out_a_valid;
	wire [2:0] domain_auto_serdesser_client_out_a_bits_opcode;
	wire [2:0] domain_auto_serdesser_client_out_a_bits_param;
	wire [3:0] domain_auto_serdesser_client_out_a_bits_size;
	wire domain_auto_serdesser_client_out_a_bits_source;
	wire [31:0] domain_auto_serdesser_client_out_a_bits_address;
	wire [3:0] domain_auto_serdesser_client_out_a_bits_mask;
	wire [31:0] domain_auto_serdesser_client_out_a_bits_data;
	wire domain_auto_serdesser_client_out_a_bits_corrupt;
	wire domain_auto_serdesser_client_out_d_ready;
	wire domain_auto_serdesser_client_out_d_valid;
	wire [2:0] domain_auto_serdesser_client_out_d_bits_opcode;
	wire [1:0] domain_auto_serdesser_client_out_d_bits_param;
	wire [3:0] domain_auto_serdesser_client_out_d_bits_size;
	wire domain_auto_serdesser_client_out_d_bits_source;
	wire domain_auto_serdesser_client_out_d_bits_sink;
	wire domain_auto_serdesser_client_out_d_bits_denied;
	wire [31:0] domain_auto_serdesser_client_out_d_bits_data;
	wire domain_auto_serdesser_client_out_d_bits_corrupt;
	wire domain_auto_tlserial_manager_crossing_in_a_ready;
	wire domain_auto_tlserial_manager_crossing_in_a_valid;
	wire [2:0] domain_auto_tlserial_manager_crossing_in_a_bits_opcode;
	wire [2:0] domain_auto_tlserial_manager_crossing_in_a_bits_param;
	wire [2:0] domain_auto_tlserial_manager_crossing_in_a_bits_size;
	wire [2:0] domain_auto_tlserial_manager_crossing_in_a_bits_source;
	wire [28:0] domain_auto_tlserial_manager_crossing_in_a_bits_address;
	wire [7:0] domain_auto_tlserial_manager_crossing_in_a_bits_mask;
	wire [63:0] domain_auto_tlserial_manager_crossing_in_a_bits_data;
	wire domain_auto_tlserial_manager_crossing_in_a_bits_corrupt;
	wire domain_auto_tlserial_manager_crossing_in_d_ready;
	wire domain_auto_tlserial_manager_crossing_in_d_valid;
	wire [2:0] domain_auto_tlserial_manager_crossing_in_d_bits_opcode;
	wire [1:0] domain_auto_tlserial_manager_crossing_in_d_bits_param;
	wire [2:0] domain_auto_tlserial_manager_crossing_in_d_bits_size;
	wire [2:0] domain_auto_tlserial_manager_crossing_in_d_bits_source;
	wire domain_auto_tlserial_manager_crossing_in_d_bits_sink;
	wire domain_auto_tlserial_manager_crossing_in_d_bits_denied;
	wire [63:0] domain_auto_tlserial_manager_crossing_in_d_bits_data;
	wire domain_auto_tlserial_manager_crossing_in_d_bits_corrupt;
	wire domain_auto_clock_in_clock;
	wire domain_auto_clock_in_reset;
	wire domain_serial_tl_in_ready;
	wire domain_serial_tl_in_valid;
	wire [31:0] domain_serial_tl_in_bits;
	wire domain_serial_tl_out_ready;
	wire domain_serial_tl_out_valid;
	wire [31:0] domain_serial_tl_out_bits;
	wire domain_clock;
	wire uartClockDomainWrapper_auto_uart_0_int_xing_out_sync_0;
	wire uartClockDomainWrapper_auto_uart_0_control_xing_in_a_ready;
	wire uartClockDomainWrapper_auto_uart_0_control_xing_in_a_valid;
	wire [2:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_opcode;
	wire [2:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_param;
	wire [1:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_size;
	wire [7:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_source;
	wire [30:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_address;
	wire [3:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_mask;
	wire [31:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_data;
	wire uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_corrupt;
	wire uartClockDomainWrapper_auto_uart_0_control_xing_in_d_ready;
	wire uartClockDomainWrapper_auto_uart_0_control_xing_in_d_valid;
	wire [2:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_opcode;
	wire [1:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_size;
	wire [7:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_source;
	wire [31:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_data;
	wire uartClockDomainWrapper_auto_uart_0_io_out_txd;
	wire uartClockDomainWrapper_auto_uart_0_io_out_rxd;
	wire uartClockDomainWrapper_auto_clock_in_clock;
	wire uartClockDomainWrapper_auto_clock_in_reset;
	wire intsink_4_auto_in_sync_0;
	wire intsink_4_auto_out_0;
	wire prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock;
	wire prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset;
	wire prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock;
	wire prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset;
	wire prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock;
	wire prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset;
	wire prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock;
	wire prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset;
	wire prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock;
	wire prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset;
	wire prci_ctrl_domain_auto_tileResetSetter_tl_in_a_ready;
	wire prci_ctrl_domain_auto_tileResetSetter_tl_in_a_valid;
	wire [2:0] prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_opcode;
	wire [2:0] prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_param;
	wire [1:0] prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_size;
	wire [7:0] prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_source;
	wire [20:0] prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_address;
	wire [3:0] prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_mask;
	wire [31:0] prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_data;
	wire prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_corrupt;
	wire prci_ctrl_domain_auto_tileResetSetter_tl_in_d_ready;
	wire prci_ctrl_domain_auto_tileResetSetter_tl_in_d_valid;
	wire [2:0] prci_ctrl_domain_auto_tileResetSetter_tl_in_d_bits_opcode;
	wire [1:0] prci_ctrl_domain_auto_tileResetSetter_tl_in_d_bits_size;
	wire [7:0] prci_ctrl_domain_auto_tileResetSetter_tl_in_d_bits_source;
	wire [31:0] prci_ctrl_domain_auto_tileResetSetter_tl_in_d_bits_data;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_ready;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_valid;
	wire [2:0] prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_opcode;
	wire [2:0] prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_param;
	wire [1:0] prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_size;
	wire [7:0] prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_source;
	wire [20:0] prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_address;
	wire [3:0] prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_mask;
	wire [31:0] prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_data;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_corrupt;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_ready;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_valid;
	wire [2:0] prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_bits_opcode;
	wire [1:0] prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_bits_size;
	wire [7:0] prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_bits_source;
	wire [31:0] prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_bits_data;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_clock;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_reset;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock;
	wire prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset;
	wire prci_ctrl_domain_auto_clock_in_clock;
	wire prci_ctrl_domain_auto_clock_in_reset;
	wire aggregator_auto_in_member_allClocks_implicit_clock_clock;
	wire aggregator_auto_in_member_allClocks_implicit_clock_reset;
	wire aggregator_auto_in_member_allClocks_subsystem_cbus_0_clock;
	wire aggregator_auto_in_member_allClocks_subsystem_cbus_0_reset;
	wire aggregator_auto_in_member_allClocks_subsystem_fbus_0_clock;
	wire aggregator_auto_in_member_allClocks_subsystem_fbus_0_reset;
	wire aggregator_auto_in_member_allClocks_subsystem_pbus_0_clock;
	wire aggregator_auto_in_member_allClocks_subsystem_pbus_0_reset;
	wire aggregator_auto_in_member_allClocks_subsystem_sbus_0_clock;
	wire aggregator_auto_in_member_allClocks_subsystem_sbus_0_reset;
	wire aggregator_auto_out_4_member_implicitClockGrouper_implicit_clock_clock;
	wire aggregator_auto_out_4_member_implicitClockGrouper_implicit_clock_reset;
	wire aggregator_auto_out_3_member_subsystem_cbus_subsystem_cbus_0_clock;
	wire aggregator_auto_out_3_member_subsystem_cbus_subsystem_cbus_0_reset;
	wire aggregator_auto_out_2_member_subsystem_fbus_subsystem_fbus_0_clock;
	wire aggregator_auto_out_2_member_subsystem_fbus_subsystem_fbus_0_reset;
	wire aggregator_auto_out_1_member_subsystem_pbus_subsystem_pbus_0_clock;
	wire aggregator_auto_out_1_member_subsystem_pbus_subsystem_pbus_0_reset;
	wire aggregator_auto_out_0_member_subsystem_sbus_subsystem_sbus_0_clock;
	wire aggregator_auto_out_0_member_subsystem_sbus_subsystem_sbus_0_reset;
	wire clockNamePrefixer_auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_clock;
	wire clockNamePrefixer_auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_reset;
	wire clockNamePrefixer_auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_clock;
	wire clockNamePrefixer_auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_reset;
	wire clockNamePrefixer_auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_clock;
	wire clockNamePrefixer_auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_reset;
	wire clockNamePrefixer_auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_clock;
	wire clockNamePrefixer_auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_reset;
	wire clockNamePrefixer_auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_clock;
	wire clockNamePrefixer_auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_reset;
	wire clockNamePrefixer_auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_clock;
	wire clockNamePrefixer_auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_reset;
	wire clockNamePrefixer_auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_clock;
	wire clockNamePrefixer_auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_reset;
	wire clockNamePrefixer_auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_clock;
	wire clockNamePrefixer_auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_reset;
	wire frequencySpecifier_auto_frequency_specifier_in_member_allClocks_implicit_clock_clock;
	wire frequencySpecifier_auto_frequency_specifier_in_member_allClocks_implicit_clock_reset;
	wire frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_clock;
	wire frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_reset;
	wire frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_clock;
	wire frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_reset;
	wire frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_clock;
	wire frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_reset;
	wire frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_clock;
	wire frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_reset;
	wire frequencySpecifier_auto_frequency_specifier_out_member_allClocks_implicit_clock_clock;
	wire frequencySpecifier_auto_frequency_specifier_out_member_allClocks_implicit_clock_reset;
	wire frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_clock;
	wire frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_reset;
	wire frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_clock;
	wire frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_reset;
	wire frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_clock;
	wire frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_reset;
	wire frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_clock;
	wire frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_reset;
	wire clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_implicit_clock_clock;
	wire clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_implicit_clock_reset;
	wire clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_clock;
	wire clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_reset;
	wire clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_clock;
	wire clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_reset;
	wire clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_clock;
	wire clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_reset;
	wire clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_clock;
	wire clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_reset;
	wire clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_implicit_clock_clock;
	wire clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_implicit_clock_reset;
	wire clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_clock;
	wire clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_reset;
	wire clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_clock;
	wire clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_reset;
	wire clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_clock;
	wire clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_reset;
	wire clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_clock;
	wire clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_reset;
	wire resetSynchronizer_auto_in_member_allClocks_implicit_clock_clock;
	wire resetSynchronizer_auto_in_member_allClocks_implicit_clock_reset;
	wire resetSynchronizer_auto_in_member_allClocks_subsystem_cbus_0_clock;
	wire resetSynchronizer_auto_in_member_allClocks_subsystem_cbus_0_reset;
	wire resetSynchronizer_auto_in_member_allClocks_subsystem_fbus_0_clock;
	wire resetSynchronizer_auto_in_member_allClocks_subsystem_fbus_0_reset;
	wire resetSynchronizer_auto_in_member_allClocks_subsystem_pbus_0_clock;
	wire resetSynchronizer_auto_in_member_allClocks_subsystem_pbus_0_reset;
	wire resetSynchronizer_auto_in_member_allClocks_subsystem_sbus_0_clock;
	wire resetSynchronizer_auto_in_member_allClocks_subsystem_sbus_0_reset;
	wire resetSynchronizer_auto_out_member_allClocks_implicit_clock_clock;
	wire resetSynchronizer_auto_out_member_allClocks_implicit_clock_reset;
	wire resetSynchronizer_auto_out_member_allClocks_subsystem_cbus_0_clock;
	wire resetSynchronizer_auto_out_member_allClocks_subsystem_cbus_0_reset;
	wire resetSynchronizer_auto_out_member_allClocks_subsystem_fbus_0_clock;
	wire resetSynchronizer_auto_out_member_allClocks_subsystem_fbus_0_reset;
	wire resetSynchronizer_auto_out_member_allClocks_subsystem_pbus_0_clock;
	wire resetSynchronizer_auto_out_member_allClocks_subsystem_pbus_0_reset;
	wire resetSynchronizer_auto_out_member_allClocks_subsystem_sbus_0_clock;
	wire resetSynchronizer_auto_out_member_allClocks_subsystem_sbus_0_reset;
	wire implicitClockGrouper_auto_in_member_implicitClockGrouper_implicit_clock_clock;
	wire implicitClockGrouper_auto_in_member_implicitClockGrouper_implicit_clock_reset;
	wire implicitClockGrouper_auto_out_clock;
	wire implicitClockGrouper_auto_out_reset;
	wire dtm_io_jtag_clock;
	wire dtm_io_jtag_reset;
	wire dtm_io_dmi_req_ready;
	wire dtm_io_dmi_req_valid;
	wire [6:0] dtm_io_dmi_req_bits_addr;
	wire [31:0] dtm_io_dmi_req_bits_data;
	wire [1:0] dtm_io_dmi_req_bits_op;
	wire dtm_io_dmi_resp_ready;
	wire dtm_io_dmi_resp_valid;
	wire [31:0] dtm_io_dmi_resp_bits_data;
	wire [1:0] dtm_io_dmi_resp_bits_resp;
	wire dtm_io_jtag_TMS;
	wire dtm_io_jtag_TDI;
	wire dtm_io_jtag_TDO_data;
	reg [6:0] int_rtc_tick_value;
	wire int_rtc_tick_wrap_wrap = int_rtc_tick_value == 7'h63;
	wire [6:0] _int_rtc_tick_wrap_value_T_1 = int_rtc_tick_value + 7'h01;
	InterruptBusWrapper ibus(
		.auto_int_bus_int_in_0(ibus_auto_int_bus_int_in_0),
		.auto_int_bus_int_out_0(ibus_auto_int_bus_int_out_0)
	);
	SystemBus subsystem_sbus(
		.auto_coupler_from_tile_tl_master_clock_xing_in_a_ready(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_ready),
		.auto_coupler_from_tile_tl_master_clock_xing_in_a_valid(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_valid),
		.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode),
		.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param),
		.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size),
		.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source),
		.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address),
		.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask),
		.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data),
		.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_corrupt(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_corrupt),
		.auto_coupler_from_tile_tl_master_clock_xing_in_d_ready(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_ready),
		.auto_coupler_from_tile_tl_master_clock_xing_in_d_valid(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_valid),
		.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode),
		.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param),
		.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size),
		.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source),
		.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink),
		.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied),
		.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data),
		.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt(subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_corrupt(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_corrupt),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data),
		.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt(subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data),
		.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt(subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt),
		.auto_fixedClockNode_out_1_clock(subsystem_sbus_auto_fixedClockNode_out_1_clock),
		.auto_fixedClockNode_out_1_reset(subsystem_sbus_auto_fixedClockNode_out_1_reset),
		.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock(subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock),
		.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset(subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset)
	);
	PeripheryBus subsystem_pbus(
		.auto_coupler_to_device_named_uart_0_control_xing_out_a_ready(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_ready),
		.auto_coupler_to_device_named_uart_0_control_xing_out_a_valid(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_valid),
		.auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode),
		.auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_param(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_param),
		.auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size),
		.auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source),
		.auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address),
		.auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask),
		.auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data),
		.auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_corrupt(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_corrupt),
		.auto_coupler_to_device_named_uart_0_control_xing_out_d_ready(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_ready),
		.auto_coupler_to_device_named_uart_0_control_xing_out_d_valid(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_valid),
		.auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode),
		.auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size),
		.auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source),
		.auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data(subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_ready(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_ready),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_valid(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_valid),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_opcode(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_opcode),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_param(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_param),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_size(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_size),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_source(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_source),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_address(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_address),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_mask(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_mask),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_data(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_data),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_corrupt(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_corrupt),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_ready(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_ready),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_valid(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_valid),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_opcode(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_opcode),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_param(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_param),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_size(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_size),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_source(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_source),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_sink(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_sink),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_denied(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_denied),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_data(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_data),
		.auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_corrupt(subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_corrupt),
		.auto_fixedClockNode_out_clock(subsystem_pbus_auto_fixedClockNode_out_clock),
		.auto_fixedClockNode_out_reset(subsystem_pbus_auto_fixedClockNode_out_reset),
		.auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock(subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock),
		.auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset(subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset),
		.auto_bus_xing_in_a_ready(subsystem_pbus_auto_bus_xing_in_a_ready),
		.auto_bus_xing_in_a_valid(subsystem_pbus_auto_bus_xing_in_a_valid),
		.auto_bus_xing_in_a_bits_opcode(subsystem_pbus_auto_bus_xing_in_a_bits_opcode),
		.auto_bus_xing_in_a_bits_param(subsystem_pbus_auto_bus_xing_in_a_bits_param),
		.auto_bus_xing_in_a_bits_size(subsystem_pbus_auto_bus_xing_in_a_bits_size),
		.auto_bus_xing_in_a_bits_source(subsystem_pbus_auto_bus_xing_in_a_bits_source),
		.auto_bus_xing_in_a_bits_address(subsystem_pbus_auto_bus_xing_in_a_bits_address),
		.auto_bus_xing_in_a_bits_mask(subsystem_pbus_auto_bus_xing_in_a_bits_mask),
		.auto_bus_xing_in_a_bits_data(subsystem_pbus_auto_bus_xing_in_a_bits_data),
		.auto_bus_xing_in_a_bits_corrupt(subsystem_pbus_auto_bus_xing_in_a_bits_corrupt),
		.auto_bus_xing_in_d_ready(subsystem_pbus_auto_bus_xing_in_d_ready),
		.auto_bus_xing_in_d_valid(subsystem_pbus_auto_bus_xing_in_d_valid),
		.auto_bus_xing_in_d_bits_opcode(subsystem_pbus_auto_bus_xing_in_d_bits_opcode),
		.auto_bus_xing_in_d_bits_param(subsystem_pbus_auto_bus_xing_in_d_bits_param),
		.auto_bus_xing_in_d_bits_size(subsystem_pbus_auto_bus_xing_in_d_bits_size),
		.auto_bus_xing_in_d_bits_source(subsystem_pbus_auto_bus_xing_in_d_bits_source),
		.auto_bus_xing_in_d_bits_sink(subsystem_pbus_auto_bus_xing_in_d_bits_sink),
		.auto_bus_xing_in_d_bits_denied(subsystem_pbus_auto_bus_xing_in_d_bits_denied),
		.auto_bus_xing_in_d_bits_data(subsystem_pbus_auto_bus_xing_in_d_bits_data),
		.auto_bus_xing_in_d_bits_corrupt(subsystem_pbus_auto_bus_xing_in_d_bits_corrupt),
		.clock(subsystem_pbus_clock),
		.reset(subsystem_pbus_reset)
	);
	FrontBus subsystem_fbus(
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_ready(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_ready),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_valid(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_valid),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_opcode(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_opcode),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_param(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_param),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_size(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_size),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_source(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_source),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_address(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_address),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_mask(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_mask),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_data(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_data),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_corrupt(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_corrupt),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_ready(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_ready),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_valid(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_valid),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_opcode(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_opcode),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_param(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_param),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_size(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_size),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_source(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_source),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_sink(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_sink),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_denied(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_denied),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_data(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_data),
		.auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_corrupt(subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_corrupt),
		.auto_fixedClockNode_out_clock(subsystem_fbus_auto_fixedClockNode_out_clock),
		.auto_fixedClockNode_out_reset(subsystem_fbus_auto_fixedClockNode_out_reset),
		.auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock(subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock),
		.auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset(subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset),
		.auto_bus_xing_out_a_ready(subsystem_fbus_auto_bus_xing_out_a_ready),
		.auto_bus_xing_out_a_valid(subsystem_fbus_auto_bus_xing_out_a_valid),
		.auto_bus_xing_out_a_bits_opcode(subsystem_fbus_auto_bus_xing_out_a_bits_opcode),
		.auto_bus_xing_out_a_bits_param(subsystem_fbus_auto_bus_xing_out_a_bits_param),
		.auto_bus_xing_out_a_bits_size(subsystem_fbus_auto_bus_xing_out_a_bits_size),
		.auto_bus_xing_out_a_bits_source(subsystem_fbus_auto_bus_xing_out_a_bits_source),
		.auto_bus_xing_out_a_bits_address(subsystem_fbus_auto_bus_xing_out_a_bits_address),
		.auto_bus_xing_out_a_bits_mask(subsystem_fbus_auto_bus_xing_out_a_bits_mask),
		.auto_bus_xing_out_a_bits_data(subsystem_fbus_auto_bus_xing_out_a_bits_data),
		.auto_bus_xing_out_a_bits_corrupt(subsystem_fbus_auto_bus_xing_out_a_bits_corrupt),
		.auto_bus_xing_out_d_ready(subsystem_fbus_auto_bus_xing_out_d_ready),
		.auto_bus_xing_out_d_valid(subsystem_fbus_auto_bus_xing_out_d_valid),
		.auto_bus_xing_out_d_bits_opcode(subsystem_fbus_auto_bus_xing_out_d_bits_opcode),
		.auto_bus_xing_out_d_bits_param(subsystem_fbus_auto_bus_xing_out_d_bits_param),
		.auto_bus_xing_out_d_bits_size(subsystem_fbus_auto_bus_xing_out_d_bits_size),
		.auto_bus_xing_out_d_bits_sink(subsystem_fbus_auto_bus_xing_out_d_bits_sink),
		.auto_bus_xing_out_d_bits_denied(subsystem_fbus_auto_bus_xing_out_d_bits_denied),
		.auto_bus_xing_out_d_bits_data(subsystem_fbus_auto_bus_xing_out_d_bits_data),
		.auto_bus_xing_out_d_bits_corrupt(subsystem_fbus_auto_bus_xing_out_d_bits_corrupt)
	);
	PeripheryBus_1 subsystem_cbus(
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_ready(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_ready),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_valid(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_valid),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_opcode(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_opcode),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_param(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_param),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_size(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_size),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_source(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_source),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_address(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_address),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_mask(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_mask),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_data(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_data),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_corrupt(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_corrupt),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_ready(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_ready),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_valid(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_valid),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_opcode(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_opcode),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_size(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_size),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_source(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_source),
		.auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_data(subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_data),
		.auto_coupler_to_slave_named_clockgater_buffer_out_a_ready(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_ready),
		.auto_coupler_to_slave_named_clockgater_buffer_out_a_valid(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_valid),
		.auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_opcode(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_opcode),
		.auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_param(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_param),
		.auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_size(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_size),
		.auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_source(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_source),
		.auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_address(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_address),
		.auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_mask(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_mask),
		.auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_data(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_data),
		.auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_corrupt(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_corrupt),
		.auto_coupler_to_slave_named_clockgater_buffer_out_d_ready(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_ready),
		.auto_coupler_to_slave_named_clockgater_buffer_out_d_valid(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_valid),
		.auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_opcode(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_opcode),
		.auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_size(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_size),
		.auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_source(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_source),
		.auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_data(subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_data),
		.auto_coupler_to_bootrom_fragmenter_out_a_ready(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_ready),
		.auto_coupler_to_bootrom_fragmenter_out_a_valid(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_valid),
		.auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode),
		.auto_coupler_to_bootrom_fragmenter_out_a_bits_param(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_param),
		.auto_coupler_to_bootrom_fragmenter_out_a_bits_size(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_size),
		.auto_coupler_to_bootrom_fragmenter_out_a_bits_source(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_source),
		.auto_coupler_to_bootrom_fragmenter_out_a_bits_address(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_address),
		.auto_coupler_to_bootrom_fragmenter_out_a_bits_mask(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_mask),
		.auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt),
		.auto_coupler_to_bootrom_fragmenter_out_d_ready(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_ready),
		.auto_coupler_to_bootrom_fragmenter_out_d_valid(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_valid),
		.auto_coupler_to_bootrom_fragmenter_out_d_bits_size(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_size),
		.auto_coupler_to_bootrom_fragmenter_out_d_bits_source(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_source),
		.auto_coupler_to_bootrom_fragmenter_out_d_bits_data(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_data),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_a_ready(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_ready),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_a_valid(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_valid),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_opcode(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_opcode),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_param(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_param),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_size(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_size),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_source(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_source),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_address(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_address),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_mask(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_mask),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_data(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_data),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_d_ready(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_ready),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_d_valid(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_valid),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_opcode(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_opcode),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_param(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_param),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_size(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_size),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_source(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_source),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_sink(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_sink),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_denied(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_denied),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_data(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_data),
		.auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_corrupt(subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_corrupt),
		.auto_coupler_to_debug_fragmenter_out_a_ready(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_ready),
		.auto_coupler_to_debug_fragmenter_out_a_valid(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_valid),
		.auto_coupler_to_debug_fragmenter_out_a_bits_opcode(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_opcode),
		.auto_coupler_to_debug_fragmenter_out_a_bits_param(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_param),
		.auto_coupler_to_debug_fragmenter_out_a_bits_size(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_size),
		.auto_coupler_to_debug_fragmenter_out_a_bits_source(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_source),
		.auto_coupler_to_debug_fragmenter_out_a_bits_address(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_address),
		.auto_coupler_to_debug_fragmenter_out_a_bits_mask(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_mask),
		.auto_coupler_to_debug_fragmenter_out_a_bits_data(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_data),
		.auto_coupler_to_debug_fragmenter_out_a_bits_corrupt(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_corrupt),
		.auto_coupler_to_debug_fragmenter_out_d_ready(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_ready),
		.auto_coupler_to_debug_fragmenter_out_d_valid(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_valid),
		.auto_coupler_to_debug_fragmenter_out_d_bits_opcode(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_bits_opcode),
		.auto_coupler_to_debug_fragmenter_out_d_bits_size(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_bits_size),
		.auto_coupler_to_debug_fragmenter_out_d_bits_source(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_bits_source),
		.auto_coupler_to_debug_fragmenter_out_d_bits_data(subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_bits_data),
		.auto_coupler_to_clint_fragmenter_out_a_ready(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_ready),
		.auto_coupler_to_clint_fragmenter_out_a_valid(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_valid),
		.auto_coupler_to_clint_fragmenter_out_a_bits_opcode(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_opcode),
		.auto_coupler_to_clint_fragmenter_out_a_bits_param(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_param),
		.auto_coupler_to_clint_fragmenter_out_a_bits_size(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_size),
		.auto_coupler_to_clint_fragmenter_out_a_bits_source(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_source),
		.auto_coupler_to_clint_fragmenter_out_a_bits_address(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_address),
		.auto_coupler_to_clint_fragmenter_out_a_bits_mask(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_mask),
		.auto_coupler_to_clint_fragmenter_out_a_bits_data(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_data),
		.auto_coupler_to_clint_fragmenter_out_a_bits_corrupt(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_corrupt),
		.auto_coupler_to_clint_fragmenter_out_d_ready(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_ready),
		.auto_coupler_to_clint_fragmenter_out_d_valid(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_valid),
		.auto_coupler_to_clint_fragmenter_out_d_bits_opcode(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_opcode),
		.auto_coupler_to_clint_fragmenter_out_d_bits_size(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_size),
		.auto_coupler_to_clint_fragmenter_out_d_bits_source(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_source),
		.auto_coupler_to_clint_fragmenter_out_d_bits_data(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_data),
		.auto_coupler_to_plic_fragmenter_out_a_ready(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_ready),
		.auto_coupler_to_plic_fragmenter_out_a_valid(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_valid),
		.auto_coupler_to_plic_fragmenter_out_a_bits_opcode(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_opcode),
		.auto_coupler_to_plic_fragmenter_out_a_bits_param(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_param),
		.auto_coupler_to_plic_fragmenter_out_a_bits_size(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_size),
		.auto_coupler_to_plic_fragmenter_out_a_bits_source(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_source),
		.auto_coupler_to_plic_fragmenter_out_a_bits_address(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_address),
		.auto_coupler_to_plic_fragmenter_out_a_bits_mask(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_mask),
		.auto_coupler_to_plic_fragmenter_out_a_bits_data(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_data),
		.auto_coupler_to_plic_fragmenter_out_a_bits_corrupt(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_corrupt),
		.auto_coupler_to_plic_fragmenter_out_d_ready(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_ready),
		.auto_coupler_to_plic_fragmenter_out_d_valid(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_valid),
		.auto_coupler_to_plic_fragmenter_out_d_bits_opcode(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_opcode),
		.auto_coupler_to_plic_fragmenter_out_d_bits_size(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_size),
		.auto_coupler_to_plic_fragmenter_out_d_bits_source(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_source),
		.auto_coupler_to_plic_fragmenter_out_d_bits_data(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_data),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_corrupt(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_corrupt),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_param(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_param),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_sink(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_sink),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data),
		.auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt(subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt),
		.auto_fixedClockNode_out_4_clock(subsystem_cbus_auto_fixedClockNode_out_4_clock),
		.auto_fixedClockNode_out_4_reset(subsystem_cbus_auto_fixedClockNode_out_4_reset),
		.auto_fixedClockNode_out_3_clock(subsystem_cbus_auto_fixedClockNode_out_3_clock),
		.auto_fixedClockNode_out_3_reset(subsystem_cbus_auto_fixedClockNode_out_3_reset),
		.auto_fixedClockNode_out_2_clock(subsystem_cbus_auto_fixedClockNode_out_2_clock),
		.auto_fixedClockNode_out_2_reset(subsystem_cbus_auto_fixedClockNode_out_2_reset),
		.auto_fixedClockNode_out_0_clock(subsystem_cbus_auto_fixedClockNode_out_0_clock),
		.auto_fixedClockNode_out_0_reset(subsystem_cbus_auto_fixedClockNode_out_0_reset),
		.auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock(subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock),
		.auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset(subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset),
		.auto_bus_xing_in_a_ready(subsystem_cbus_auto_bus_xing_in_a_ready),
		.auto_bus_xing_in_a_valid(subsystem_cbus_auto_bus_xing_in_a_valid),
		.auto_bus_xing_in_a_bits_opcode(subsystem_cbus_auto_bus_xing_in_a_bits_opcode),
		.auto_bus_xing_in_a_bits_param(subsystem_cbus_auto_bus_xing_in_a_bits_param),
		.auto_bus_xing_in_a_bits_size(subsystem_cbus_auto_bus_xing_in_a_bits_size),
		.auto_bus_xing_in_a_bits_source(subsystem_cbus_auto_bus_xing_in_a_bits_source),
		.auto_bus_xing_in_a_bits_address(subsystem_cbus_auto_bus_xing_in_a_bits_address),
		.auto_bus_xing_in_a_bits_mask(subsystem_cbus_auto_bus_xing_in_a_bits_mask),
		.auto_bus_xing_in_a_bits_data(subsystem_cbus_auto_bus_xing_in_a_bits_data),
		.auto_bus_xing_in_a_bits_corrupt(subsystem_cbus_auto_bus_xing_in_a_bits_corrupt),
		.auto_bus_xing_in_d_ready(subsystem_cbus_auto_bus_xing_in_d_ready),
		.auto_bus_xing_in_d_valid(subsystem_cbus_auto_bus_xing_in_d_valid),
		.auto_bus_xing_in_d_bits_opcode(subsystem_cbus_auto_bus_xing_in_d_bits_opcode),
		.auto_bus_xing_in_d_bits_param(subsystem_cbus_auto_bus_xing_in_d_bits_param),
		.auto_bus_xing_in_d_bits_size(subsystem_cbus_auto_bus_xing_in_d_bits_size),
		.auto_bus_xing_in_d_bits_source(subsystem_cbus_auto_bus_xing_in_d_bits_source),
		.auto_bus_xing_in_d_bits_sink(subsystem_cbus_auto_bus_xing_in_d_bits_sink),
		.auto_bus_xing_in_d_bits_denied(subsystem_cbus_auto_bus_xing_in_d_bits_denied),
		.auto_bus_xing_in_d_bits_data(subsystem_cbus_auto_bus_xing_in_d_bits_data),
		.auto_bus_xing_in_d_bits_corrupt(subsystem_cbus_auto_bus_xing_in_d_bits_corrupt),
		.custom_boot(subsystem_cbus_custom_boot),
		.clock(subsystem_cbus_clock),
		.reset(subsystem_cbus_reset)
	);
	TilePRCIDomain tile_prci_domain(
		.auto_intsink_in_sync_0(tile_prci_domain_auto_intsink_in_sync_0),
		.auto_tile_reset_domain_tile_hartid_in(tile_prci_domain_auto_tile_reset_domain_tile_hartid_in),
		.auto_int_out_clock_xing_out_2_sync_0(tile_prci_domain_auto_int_out_clock_xing_out_2_sync_0),
		.auto_int_out_clock_xing_out_1_sync_0(tile_prci_domain_auto_int_out_clock_xing_out_1_sync_0),
		.auto_int_out_clock_xing_out_0_sync_0(tile_prci_domain_auto_int_out_clock_xing_out_0_sync_0),
		.auto_int_in_clock_xing_in_1_sync_0(tile_prci_domain_auto_int_in_clock_xing_in_1_sync_0),
		.auto_int_in_clock_xing_in_0_sync_0(tile_prci_domain_auto_int_in_clock_xing_in_0_sync_0),
		.auto_int_in_clock_xing_in_0_sync_1(tile_prci_domain_auto_int_in_clock_xing_in_0_sync_1),
		.auto_tl_slave_clock_xing_in_a_ready(tile_prci_domain_auto_tl_slave_clock_xing_in_a_ready),
		.auto_tl_slave_clock_xing_in_a_valid(tile_prci_domain_auto_tl_slave_clock_xing_in_a_valid),
		.auto_tl_slave_clock_xing_in_a_bits_opcode(tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_opcode),
		.auto_tl_slave_clock_xing_in_a_bits_param(tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_param),
		.auto_tl_slave_clock_xing_in_a_bits_size(tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_size),
		.auto_tl_slave_clock_xing_in_a_bits_source(tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_source),
		.auto_tl_slave_clock_xing_in_a_bits_address(tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_address),
		.auto_tl_slave_clock_xing_in_a_bits_mask(tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_mask),
		.auto_tl_slave_clock_xing_in_a_bits_data(tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_data),
		.auto_tl_slave_clock_xing_in_d_ready(tile_prci_domain_auto_tl_slave_clock_xing_in_d_ready),
		.auto_tl_slave_clock_xing_in_d_valid(tile_prci_domain_auto_tl_slave_clock_xing_in_d_valid),
		.auto_tl_slave_clock_xing_in_d_bits_opcode(tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_opcode),
		.auto_tl_slave_clock_xing_in_d_bits_param(tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_param),
		.auto_tl_slave_clock_xing_in_d_bits_size(tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_size),
		.auto_tl_slave_clock_xing_in_d_bits_source(tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_source),
		.auto_tl_slave_clock_xing_in_d_bits_sink(tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_sink),
		.auto_tl_slave_clock_xing_in_d_bits_denied(tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_denied),
		.auto_tl_slave_clock_xing_in_d_bits_data(tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_data),
		.auto_tl_slave_clock_xing_in_d_bits_corrupt(tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_corrupt),
		.auto_tl_master_clock_xing_out_a_ready(tile_prci_domain_auto_tl_master_clock_xing_out_a_ready),
		.auto_tl_master_clock_xing_out_a_valid(tile_prci_domain_auto_tl_master_clock_xing_out_a_valid),
		.auto_tl_master_clock_xing_out_a_bits_opcode(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_opcode),
		.auto_tl_master_clock_xing_out_a_bits_param(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_param),
		.auto_tl_master_clock_xing_out_a_bits_size(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_size),
		.auto_tl_master_clock_xing_out_a_bits_source(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_source),
		.auto_tl_master_clock_xing_out_a_bits_address(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_address),
		.auto_tl_master_clock_xing_out_a_bits_mask(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_mask),
		.auto_tl_master_clock_xing_out_a_bits_data(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_data),
		.auto_tl_master_clock_xing_out_a_bits_corrupt(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_corrupt),
		.auto_tl_master_clock_xing_out_d_ready(tile_prci_domain_auto_tl_master_clock_xing_out_d_ready),
		.auto_tl_master_clock_xing_out_d_valid(tile_prci_domain_auto_tl_master_clock_xing_out_d_valid),
		.auto_tl_master_clock_xing_out_d_bits_opcode(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_opcode),
		.auto_tl_master_clock_xing_out_d_bits_param(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_param),
		.auto_tl_master_clock_xing_out_d_bits_size(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_size),
		.auto_tl_master_clock_xing_out_d_bits_source(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_source),
		.auto_tl_master_clock_xing_out_d_bits_sink(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_sink),
		.auto_tl_master_clock_xing_out_d_bits_denied(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_denied),
		.auto_tl_master_clock_xing_out_d_bits_data(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_data),
		.auto_tl_master_clock_xing_out_d_bits_corrupt(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_corrupt),
		.auto_tap_clock_in_clock(tile_prci_domain_auto_tap_clock_in_clock),
		.auto_tap_clock_in_reset(tile_prci_domain_auto_tap_clock_in_reset)
	);
	ClockSinkDomain plicDomainWrapper(
		.auto_plic_int_in_0(plicDomainWrapper_auto_plic_int_in_0),
		.auto_plic_int_out_0(plicDomainWrapper_auto_plic_int_out_0),
		.auto_plic_in_a_ready(plicDomainWrapper_auto_plic_in_a_ready),
		.auto_plic_in_a_valid(plicDomainWrapper_auto_plic_in_a_valid),
		.auto_plic_in_a_bits_opcode(plicDomainWrapper_auto_plic_in_a_bits_opcode),
		.auto_plic_in_a_bits_param(plicDomainWrapper_auto_plic_in_a_bits_param),
		.auto_plic_in_a_bits_size(plicDomainWrapper_auto_plic_in_a_bits_size),
		.auto_plic_in_a_bits_source(plicDomainWrapper_auto_plic_in_a_bits_source),
		.auto_plic_in_a_bits_address(plicDomainWrapper_auto_plic_in_a_bits_address),
		.auto_plic_in_a_bits_mask(plicDomainWrapper_auto_plic_in_a_bits_mask),
		.auto_plic_in_a_bits_data(plicDomainWrapper_auto_plic_in_a_bits_data),
		.auto_plic_in_a_bits_corrupt(plicDomainWrapper_auto_plic_in_a_bits_corrupt),
		.auto_plic_in_d_ready(plicDomainWrapper_auto_plic_in_d_ready),
		.auto_plic_in_d_valid(plicDomainWrapper_auto_plic_in_d_valid),
		.auto_plic_in_d_bits_opcode(plicDomainWrapper_auto_plic_in_d_bits_opcode),
		.auto_plic_in_d_bits_size(plicDomainWrapper_auto_plic_in_d_bits_size),
		.auto_plic_in_d_bits_source(plicDomainWrapper_auto_plic_in_d_bits_source),
		.auto_plic_in_d_bits_data(plicDomainWrapper_auto_plic_in_d_bits_data),
		.auto_clock_in_clock(plicDomainWrapper_auto_clock_in_clock),
		.auto_clock_in_reset(plicDomainWrapper_auto_clock_in_reset)
	);
	CLINT clint(
		.clock(clint_clock),
		.reset(clint_reset),
		.auto_int_out_0(clint_auto_int_out_0),
		.auto_int_out_1(clint_auto_int_out_1),
		.auto_in_a_ready(clint_auto_in_a_ready),
		.auto_in_a_valid(clint_auto_in_a_valid),
		.auto_in_a_bits_opcode(clint_auto_in_a_bits_opcode),
		.auto_in_a_bits_param(clint_auto_in_a_bits_param),
		.auto_in_a_bits_size(clint_auto_in_a_bits_size),
		.auto_in_a_bits_source(clint_auto_in_a_bits_source),
		.auto_in_a_bits_address(clint_auto_in_a_bits_address),
		.auto_in_a_bits_mask(clint_auto_in_a_bits_mask),
		.auto_in_a_bits_data(clint_auto_in_a_bits_data),
		.auto_in_a_bits_corrupt(clint_auto_in_a_bits_corrupt),
		.auto_in_d_ready(clint_auto_in_d_ready),
		.auto_in_d_valid(clint_auto_in_d_valid),
		.auto_in_d_bits_opcode(clint_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(clint_auto_in_d_bits_size),
		.auto_in_d_bits_source(clint_auto_in_d_bits_source),
		.auto_in_d_bits_data(clint_auto_in_d_bits_data),
		.io_rtcTick(clint_io_rtcTick)
	);
	TLDebugModule debug_1(
		.auto_dmInner_dmInner_tl_in_a_ready(debug_1_auto_dmInner_dmInner_tl_in_a_ready),
		.auto_dmInner_dmInner_tl_in_a_valid(debug_1_auto_dmInner_dmInner_tl_in_a_valid),
		.auto_dmInner_dmInner_tl_in_a_bits_opcode(debug_1_auto_dmInner_dmInner_tl_in_a_bits_opcode),
		.auto_dmInner_dmInner_tl_in_a_bits_param(debug_1_auto_dmInner_dmInner_tl_in_a_bits_param),
		.auto_dmInner_dmInner_tl_in_a_bits_size(debug_1_auto_dmInner_dmInner_tl_in_a_bits_size),
		.auto_dmInner_dmInner_tl_in_a_bits_source(debug_1_auto_dmInner_dmInner_tl_in_a_bits_source),
		.auto_dmInner_dmInner_tl_in_a_bits_address(debug_1_auto_dmInner_dmInner_tl_in_a_bits_address),
		.auto_dmInner_dmInner_tl_in_a_bits_mask(debug_1_auto_dmInner_dmInner_tl_in_a_bits_mask),
		.auto_dmInner_dmInner_tl_in_a_bits_data(debug_1_auto_dmInner_dmInner_tl_in_a_bits_data),
		.auto_dmInner_dmInner_tl_in_a_bits_corrupt(debug_1_auto_dmInner_dmInner_tl_in_a_bits_corrupt),
		.auto_dmInner_dmInner_tl_in_d_ready(debug_1_auto_dmInner_dmInner_tl_in_d_ready),
		.auto_dmInner_dmInner_tl_in_d_valid(debug_1_auto_dmInner_dmInner_tl_in_d_valid),
		.auto_dmInner_dmInner_tl_in_d_bits_opcode(debug_1_auto_dmInner_dmInner_tl_in_d_bits_opcode),
		.auto_dmInner_dmInner_tl_in_d_bits_size(debug_1_auto_dmInner_dmInner_tl_in_d_bits_size),
		.auto_dmInner_dmInner_tl_in_d_bits_source(debug_1_auto_dmInner_dmInner_tl_in_d_bits_source),
		.auto_dmInner_dmInner_tl_in_d_bits_data(debug_1_auto_dmInner_dmInner_tl_in_d_bits_data),
		.auto_dmOuter_intsource_out_sync_0(debug_1_auto_dmOuter_intsource_out_sync_0),
		.io_debug_clock(debug_1_io_debug_clock),
		.io_debug_reset(debug_1_io_debug_reset),
		.io_ctrl_dmactive(debug_1_io_ctrl_dmactive),
		.io_ctrl_dmactiveAck(debug_1_io_ctrl_dmactiveAck),
		.io_dmi_dmi_req_ready(debug_1_io_dmi_dmi_req_ready),
		.io_dmi_dmi_req_valid(debug_1_io_dmi_dmi_req_valid),
		.io_dmi_dmi_req_bits_addr(debug_1_io_dmi_dmi_req_bits_addr),
		.io_dmi_dmi_req_bits_data(debug_1_io_dmi_dmi_req_bits_data),
		.io_dmi_dmi_req_bits_op(debug_1_io_dmi_dmi_req_bits_op),
		.io_dmi_dmi_resp_ready(debug_1_io_dmi_dmi_resp_ready),
		.io_dmi_dmi_resp_valid(debug_1_io_dmi_dmi_resp_valid),
		.io_dmi_dmi_resp_bits_data(debug_1_io_dmi_dmi_resp_bits_data),
		.io_dmi_dmi_resp_bits_resp(debug_1_io_dmi_dmi_resp_bits_resp),
		.io_dmi_dmiClock(debug_1_io_dmi_dmiClock),
		.io_dmi_dmiReset(debug_1_io_dmi_dmiReset),
		.io_hartIsInReset_0(debug_1_io_hartIsInReset_0)
	);
	IntXbar xbar(
		.auto_int_in_0(xbar_auto_int_in_0),
		.auto_int_out_0(xbar_auto_int_out_0)
	);
	IntXbar xbar_1(
		.auto_int_in_0(xbar_1_auto_int_in_0),
		.auto_int_out_0(xbar_1_auto_int_out_0)
	);
	IntXbar xbar_2(
		.auto_int_in_0(xbar_2_auto_int_in_0),
		.auto_int_out_0(xbar_2_auto_int_out_0)
	);
	BundleBridgeNexus_13 tileHartIdNexusNode(.auto_out(tileHartIdNexusNode_auto_out));
	IntSyncCrossingSource_5 intsource(
		.clock(intsource_clock),
		.reset(intsource_reset),
		.auto_in_0(intsource_auto_in_0),
		.auto_in_1(intsource_auto_in_1),
		.auto_out_sync_0(intsource_auto_out_sync_0),
		.auto_out_sync_1(intsource_auto_out_sync_1)
	);
	IntSyncCrossingSource_1 intsource_1(
		.clock(intsource_1_clock),
		.reset(intsource_1_reset),
		.auto_in_0(intsource_1_auto_in_0),
		.auto_out_sync_0(intsource_1_auto_out_sync_0)
	);
	IntSyncSyncCrossingSink_1 intsink_1(
		.auto_in_sync_0(intsink_1_auto_in_sync_0),
		.auto_out_0(intsink_1_auto_out_0)
	);
	IntSyncSyncCrossingSink_1 intsink_2(
		.auto_in_sync_0(intsink_2_auto_in_sync_0),
		.auto_out_0(intsink_2_auto_out_0)
	);
	IntSyncSyncCrossingSink_1 intsink_3(
		.auto_in_sync_0(intsink_3_auto_in_sync_0),
		.auto_out_0(intsink_3_auto_out_0)
	);
	ClockSinkDomain_1 bootROMDomainWrapper(
		.auto_bootrom_in_a_ready(bootROMDomainWrapper_auto_bootrom_in_a_ready),
		.auto_bootrom_in_a_valid(bootROMDomainWrapper_auto_bootrom_in_a_valid),
		.auto_bootrom_in_a_bits_opcode(bootROMDomainWrapper_auto_bootrom_in_a_bits_opcode),
		.auto_bootrom_in_a_bits_param(bootROMDomainWrapper_auto_bootrom_in_a_bits_param),
		.auto_bootrom_in_a_bits_size(bootROMDomainWrapper_auto_bootrom_in_a_bits_size),
		.auto_bootrom_in_a_bits_source(bootROMDomainWrapper_auto_bootrom_in_a_bits_source),
		.auto_bootrom_in_a_bits_address(bootROMDomainWrapper_auto_bootrom_in_a_bits_address),
		.auto_bootrom_in_a_bits_mask(bootROMDomainWrapper_auto_bootrom_in_a_bits_mask),
		.auto_bootrom_in_a_bits_corrupt(bootROMDomainWrapper_auto_bootrom_in_a_bits_corrupt),
		.auto_bootrom_in_d_ready(bootROMDomainWrapper_auto_bootrom_in_d_ready),
		.auto_bootrom_in_d_valid(bootROMDomainWrapper_auto_bootrom_in_d_valid),
		.auto_bootrom_in_d_bits_size(bootROMDomainWrapper_auto_bootrom_in_d_bits_size),
		.auto_bootrom_in_d_bits_source(bootROMDomainWrapper_auto_bootrom_in_d_bits_source),
		.auto_bootrom_in_d_bits_data(bootROMDomainWrapper_auto_bootrom_in_d_bits_data),
		.auto_clock_in_clock(bootROMDomainWrapper_auto_clock_in_clock),
		.auto_clock_in_reset(bootROMDomainWrapper_auto_clock_in_reset)
	);
	ClockSinkDomain_2 domain(
		.auto_serdesser_client_out_a_ready(domain_auto_serdesser_client_out_a_ready),
		.auto_serdesser_client_out_a_valid(domain_auto_serdesser_client_out_a_valid),
		.auto_serdesser_client_out_a_bits_opcode(domain_auto_serdesser_client_out_a_bits_opcode),
		.auto_serdesser_client_out_a_bits_param(domain_auto_serdesser_client_out_a_bits_param),
		.auto_serdesser_client_out_a_bits_size(domain_auto_serdesser_client_out_a_bits_size),
		.auto_serdesser_client_out_a_bits_source(domain_auto_serdesser_client_out_a_bits_source),
		.auto_serdesser_client_out_a_bits_address(domain_auto_serdesser_client_out_a_bits_address),
		.auto_serdesser_client_out_a_bits_mask(domain_auto_serdesser_client_out_a_bits_mask),
		.auto_serdesser_client_out_a_bits_data(domain_auto_serdesser_client_out_a_bits_data),
		.auto_serdesser_client_out_a_bits_corrupt(domain_auto_serdesser_client_out_a_bits_corrupt),
		.auto_serdesser_client_out_d_ready(domain_auto_serdesser_client_out_d_ready),
		.auto_serdesser_client_out_d_valid(domain_auto_serdesser_client_out_d_valid),
		.auto_serdesser_client_out_d_bits_opcode(domain_auto_serdesser_client_out_d_bits_opcode),
		.auto_serdesser_client_out_d_bits_param(domain_auto_serdesser_client_out_d_bits_param),
		.auto_serdesser_client_out_d_bits_size(domain_auto_serdesser_client_out_d_bits_size),
		.auto_serdesser_client_out_d_bits_source(domain_auto_serdesser_client_out_d_bits_source),
		.auto_serdesser_client_out_d_bits_sink(domain_auto_serdesser_client_out_d_bits_sink),
		.auto_serdesser_client_out_d_bits_denied(domain_auto_serdesser_client_out_d_bits_denied),
		.auto_serdesser_client_out_d_bits_data(domain_auto_serdesser_client_out_d_bits_data),
		.auto_serdesser_client_out_d_bits_corrupt(domain_auto_serdesser_client_out_d_bits_corrupt),
		.auto_tlserial_manager_crossing_in_a_ready(domain_auto_tlserial_manager_crossing_in_a_ready),
		.auto_tlserial_manager_crossing_in_a_valid(domain_auto_tlserial_manager_crossing_in_a_valid),
		.auto_tlserial_manager_crossing_in_a_bits_opcode(domain_auto_tlserial_manager_crossing_in_a_bits_opcode),
		.auto_tlserial_manager_crossing_in_a_bits_param(domain_auto_tlserial_manager_crossing_in_a_bits_param),
		.auto_tlserial_manager_crossing_in_a_bits_size(domain_auto_tlserial_manager_crossing_in_a_bits_size),
		.auto_tlserial_manager_crossing_in_a_bits_source(domain_auto_tlserial_manager_crossing_in_a_bits_source),
		.auto_tlserial_manager_crossing_in_a_bits_address(domain_auto_tlserial_manager_crossing_in_a_bits_address),
		.auto_tlserial_manager_crossing_in_a_bits_mask(domain_auto_tlserial_manager_crossing_in_a_bits_mask),
		.auto_tlserial_manager_crossing_in_a_bits_data(domain_auto_tlserial_manager_crossing_in_a_bits_data),
		.auto_tlserial_manager_crossing_in_a_bits_corrupt(domain_auto_tlserial_manager_crossing_in_a_bits_corrupt),
		.auto_tlserial_manager_crossing_in_d_ready(domain_auto_tlserial_manager_crossing_in_d_ready),
		.auto_tlserial_manager_crossing_in_d_valid(domain_auto_tlserial_manager_crossing_in_d_valid),
		.auto_tlserial_manager_crossing_in_d_bits_opcode(domain_auto_tlserial_manager_crossing_in_d_bits_opcode),
		.auto_tlserial_manager_crossing_in_d_bits_param(domain_auto_tlserial_manager_crossing_in_d_bits_param),
		.auto_tlserial_manager_crossing_in_d_bits_size(domain_auto_tlserial_manager_crossing_in_d_bits_size),
		.auto_tlserial_manager_crossing_in_d_bits_source(domain_auto_tlserial_manager_crossing_in_d_bits_source),
		.auto_tlserial_manager_crossing_in_d_bits_sink(domain_auto_tlserial_manager_crossing_in_d_bits_sink),
		.auto_tlserial_manager_crossing_in_d_bits_denied(domain_auto_tlserial_manager_crossing_in_d_bits_denied),
		.auto_tlserial_manager_crossing_in_d_bits_data(domain_auto_tlserial_manager_crossing_in_d_bits_data),
		.auto_tlserial_manager_crossing_in_d_bits_corrupt(domain_auto_tlserial_manager_crossing_in_d_bits_corrupt),
		.auto_clock_in_clock(domain_auto_clock_in_clock),
		.auto_clock_in_reset(domain_auto_clock_in_reset),
		.serial_tl_in_ready(domain_serial_tl_in_ready),
		.serial_tl_in_valid(domain_serial_tl_in_valid),
		.serial_tl_in_bits(domain_serial_tl_in_bits),
		.serial_tl_out_ready(domain_serial_tl_out_ready),
		.serial_tl_out_valid(domain_serial_tl_out_valid),
		.serial_tl_out_bits(domain_serial_tl_out_bits),
		.clock(domain_clock)
	);
	ClockSinkDomain_3 uartClockDomainWrapper(
		.auto_uart_0_int_xing_out_sync_0(uartClockDomainWrapper_auto_uart_0_int_xing_out_sync_0),
		.auto_uart_0_control_xing_in_a_ready(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_ready),
		.auto_uart_0_control_xing_in_a_valid(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_valid),
		.auto_uart_0_control_xing_in_a_bits_opcode(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_opcode),
		.auto_uart_0_control_xing_in_a_bits_param(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_param),
		.auto_uart_0_control_xing_in_a_bits_size(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_size),
		.auto_uart_0_control_xing_in_a_bits_source(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_source),
		.auto_uart_0_control_xing_in_a_bits_address(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_address),
		.auto_uart_0_control_xing_in_a_bits_mask(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_mask),
		.auto_uart_0_control_xing_in_a_bits_data(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_data),
		.auto_uart_0_control_xing_in_a_bits_corrupt(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_corrupt),
		.auto_uart_0_control_xing_in_d_ready(uartClockDomainWrapper_auto_uart_0_control_xing_in_d_ready),
		.auto_uart_0_control_xing_in_d_valid(uartClockDomainWrapper_auto_uart_0_control_xing_in_d_valid),
		.auto_uart_0_control_xing_in_d_bits_opcode(uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_opcode),
		.auto_uart_0_control_xing_in_d_bits_size(uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_size),
		.auto_uart_0_control_xing_in_d_bits_source(uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_source),
		.auto_uart_0_control_xing_in_d_bits_data(uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_data),
		.auto_uart_0_io_out_txd(uartClockDomainWrapper_auto_uart_0_io_out_txd),
		.auto_uart_0_io_out_rxd(uartClockDomainWrapper_auto_uart_0_io_out_rxd),
		.auto_clock_in_clock(uartClockDomainWrapper_auto_clock_in_clock),
		.auto_clock_in_reset(uartClockDomainWrapper_auto_clock_in_reset)
	);
	IntSyncSyncCrossingSink_1 intsink_4(
		.auto_in_sync_0(intsink_4_auto_in_sync_0),
		.auto_out_0(intsink_4_auto_out_0)
	);
	ClockSinkDomain_4 prci_ctrl_domain(
		.auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock(prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock),
		.auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset(prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset),
		.auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock(prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock),
		.auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset(prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset),
		.auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock(prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock),
		.auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset(prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset),
		.auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock(prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock),
		.auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset(prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset),
		.auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock(prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock),
		.auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset(prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset),
		.auto_tileResetSetter_tl_in_a_ready(prci_ctrl_domain_auto_tileResetSetter_tl_in_a_ready),
		.auto_tileResetSetter_tl_in_a_valid(prci_ctrl_domain_auto_tileResetSetter_tl_in_a_valid),
		.auto_tileResetSetter_tl_in_a_bits_opcode(prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_opcode),
		.auto_tileResetSetter_tl_in_a_bits_param(prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_param),
		.auto_tileResetSetter_tl_in_a_bits_size(prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_size),
		.auto_tileResetSetter_tl_in_a_bits_source(prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_source),
		.auto_tileResetSetter_tl_in_a_bits_address(prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_address),
		.auto_tileResetSetter_tl_in_a_bits_mask(prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_mask),
		.auto_tileResetSetter_tl_in_a_bits_data(prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_data),
		.auto_tileResetSetter_tl_in_a_bits_corrupt(prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_corrupt),
		.auto_tileResetSetter_tl_in_d_ready(prci_ctrl_domain_auto_tileResetSetter_tl_in_d_ready),
		.auto_tileResetSetter_tl_in_d_valid(prci_ctrl_domain_auto_tileResetSetter_tl_in_d_valid),
		.auto_tileResetSetter_tl_in_d_bits_opcode(prci_ctrl_domain_auto_tileResetSetter_tl_in_d_bits_opcode),
		.auto_tileResetSetter_tl_in_d_bits_size(prci_ctrl_domain_auto_tileResetSetter_tl_in_d_bits_size),
		.auto_tileResetSetter_tl_in_d_bits_source(prci_ctrl_domain_auto_tileResetSetter_tl_in_d_bits_source),
		.auto_tileResetSetter_tl_in_d_bits_data(prci_ctrl_domain_auto_tileResetSetter_tl_in_d_bits_data),
		.auto_tileClockGater_tile_clock_gater_in_a_ready(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_ready),
		.auto_tileClockGater_tile_clock_gater_in_a_valid(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_valid),
		.auto_tileClockGater_tile_clock_gater_in_a_bits_opcode(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_opcode),
		.auto_tileClockGater_tile_clock_gater_in_a_bits_param(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_param),
		.auto_tileClockGater_tile_clock_gater_in_a_bits_size(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_size),
		.auto_tileClockGater_tile_clock_gater_in_a_bits_source(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_source),
		.auto_tileClockGater_tile_clock_gater_in_a_bits_address(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_address),
		.auto_tileClockGater_tile_clock_gater_in_a_bits_mask(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_mask),
		.auto_tileClockGater_tile_clock_gater_in_a_bits_data(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_data),
		.auto_tileClockGater_tile_clock_gater_in_a_bits_corrupt(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_corrupt),
		.auto_tileClockGater_tile_clock_gater_in_d_ready(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_ready),
		.auto_tileClockGater_tile_clock_gater_in_d_valid(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_valid),
		.auto_tileClockGater_tile_clock_gater_in_d_bits_opcode(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_bits_opcode),
		.auto_tileClockGater_tile_clock_gater_in_d_bits_size(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_bits_size),
		.auto_tileClockGater_tile_clock_gater_in_d_bits_source(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_bits_source),
		.auto_tileClockGater_tile_clock_gater_in_d_bits_data(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_bits_data),
		.auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_clock(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_clock),
		.auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_reset(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_reset),
		.auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock),
		.auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset),
		.auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock),
		.auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset),
		.auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock),
		.auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset),
		.auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock),
		.auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset(prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset),
		.auto_clock_in_clock(prci_ctrl_domain_auto_clock_in_clock),
		.auto_clock_in_reset(prci_ctrl_domain_auto_clock_in_reset)
	);
	ClockGroupAggregator_4 aggregator(
		.auto_in_member_allClocks_implicit_clock_clock(aggregator_auto_in_member_allClocks_implicit_clock_clock),
		.auto_in_member_allClocks_implicit_clock_reset(aggregator_auto_in_member_allClocks_implicit_clock_reset),
		.auto_in_member_allClocks_subsystem_cbus_0_clock(aggregator_auto_in_member_allClocks_subsystem_cbus_0_clock),
		.auto_in_member_allClocks_subsystem_cbus_0_reset(aggregator_auto_in_member_allClocks_subsystem_cbus_0_reset),
		.auto_in_member_allClocks_subsystem_fbus_0_clock(aggregator_auto_in_member_allClocks_subsystem_fbus_0_clock),
		.auto_in_member_allClocks_subsystem_fbus_0_reset(aggregator_auto_in_member_allClocks_subsystem_fbus_0_reset),
		.auto_in_member_allClocks_subsystem_pbus_0_clock(aggregator_auto_in_member_allClocks_subsystem_pbus_0_clock),
		.auto_in_member_allClocks_subsystem_pbus_0_reset(aggregator_auto_in_member_allClocks_subsystem_pbus_0_reset),
		.auto_in_member_allClocks_subsystem_sbus_0_clock(aggregator_auto_in_member_allClocks_subsystem_sbus_0_clock),
		.auto_in_member_allClocks_subsystem_sbus_0_reset(aggregator_auto_in_member_allClocks_subsystem_sbus_0_reset),
		.auto_out_4_member_implicitClockGrouper_implicit_clock_clock(aggregator_auto_out_4_member_implicitClockGrouper_implicit_clock_clock),
		.auto_out_4_member_implicitClockGrouper_implicit_clock_reset(aggregator_auto_out_4_member_implicitClockGrouper_implicit_clock_reset),
		.auto_out_3_member_subsystem_cbus_subsystem_cbus_0_clock(aggregator_auto_out_3_member_subsystem_cbus_subsystem_cbus_0_clock),
		.auto_out_3_member_subsystem_cbus_subsystem_cbus_0_reset(aggregator_auto_out_3_member_subsystem_cbus_subsystem_cbus_0_reset),
		.auto_out_2_member_subsystem_fbus_subsystem_fbus_0_clock(aggregator_auto_out_2_member_subsystem_fbus_subsystem_fbus_0_clock),
		.auto_out_2_member_subsystem_fbus_subsystem_fbus_0_reset(aggregator_auto_out_2_member_subsystem_fbus_subsystem_fbus_0_reset),
		.auto_out_1_member_subsystem_pbus_subsystem_pbus_0_clock(aggregator_auto_out_1_member_subsystem_pbus_subsystem_pbus_0_clock),
		.auto_out_1_member_subsystem_pbus_subsystem_pbus_0_reset(aggregator_auto_out_1_member_subsystem_pbus_subsystem_pbus_0_reset),
		.auto_out_0_member_subsystem_sbus_subsystem_sbus_0_clock(aggregator_auto_out_0_member_subsystem_sbus_subsystem_sbus_0_clock),
		.auto_out_0_member_subsystem_sbus_subsystem_sbus_0_reset(aggregator_auto_out_0_member_subsystem_sbus_subsystem_sbus_0_reset)
	);
	ClockGroupParameterModifier clockNamePrefixer(
		.auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_clock(clockNamePrefixer_auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_clock),
		.auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_reset(clockNamePrefixer_auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_reset),
		.auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_clock(clockNamePrefixer_auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_clock),
		.auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_reset(clockNamePrefixer_auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_reset),
		.auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_clock(clockNamePrefixer_auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_clock),
		.auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_reset(clockNamePrefixer_auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_reset),
		.auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_clock(clockNamePrefixer_auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_clock),
		.auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_reset(clockNamePrefixer_auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_reset),
		.auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_clock(clockNamePrefixer_auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_clock),
		.auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_reset(clockNamePrefixer_auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_reset),
		.auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_clock(clockNamePrefixer_auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_clock),
		.auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_reset(clockNamePrefixer_auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_reset),
		.auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_clock(clockNamePrefixer_auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_clock),
		.auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_reset(clockNamePrefixer_auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_reset),
		.auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_clock(clockNamePrefixer_auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_clock),
		.auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_reset(clockNamePrefixer_auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_reset)
	);
	ClockGroupParameterModifier_1 frequencySpecifier(
		.auto_frequency_specifier_in_member_allClocks_implicit_clock_clock(frequencySpecifier_auto_frequency_specifier_in_member_allClocks_implicit_clock_clock),
		.auto_frequency_specifier_in_member_allClocks_implicit_clock_reset(frequencySpecifier_auto_frequency_specifier_in_member_allClocks_implicit_clock_reset),
		.auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_clock(frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_clock),
		.auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_reset(frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_reset),
		.auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_clock(frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_clock),
		.auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_reset(frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_reset),
		.auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_clock(frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_clock),
		.auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_reset(frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_reset),
		.auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_clock(frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_clock),
		.auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_reset(frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_reset),
		.auto_frequency_specifier_out_member_allClocks_implicit_clock_clock(frequencySpecifier_auto_frequency_specifier_out_member_allClocks_implicit_clock_clock),
		.auto_frequency_specifier_out_member_allClocks_implicit_clock_reset(frequencySpecifier_auto_frequency_specifier_out_member_allClocks_implicit_clock_reset),
		.auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_clock(frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_clock),
		.auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_reset(frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_reset),
		.auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_clock(frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_clock),
		.auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_reset(frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_reset),
		.auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_clock(frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_clock),
		.auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_reset(frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_reset),
		.auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_clock(frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_clock),
		.auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_reset(frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_reset)
	);
	ClockGroupCombiner clockGroupCombiner(
		.auto_clock_group_combiner_in_member_allClocks_implicit_clock_clock(clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_implicit_clock_clock),
		.auto_clock_group_combiner_in_member_allClocks_implicit_clock_reset(clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_implicit_clock_reset),
		.auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_clock(clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_clock),
		.auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_reset(clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_reset),
		.auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_clock(clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_clock),
		.auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_reset(clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_reset),
		.auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_clock(clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_clock),
		.auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_reset(clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_reset),
		.auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_clock(clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_clock),
		.auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_reset(clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_reset),
		.auto_clock_group_combiner_out_member_allClocks_implicit_clock_clock(clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_implicit_clock_clock),
		.auto_clock_group_combiner_out_member_allClocks_implicit_clock_reset(clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_implicit_clock_reset),
		.auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_clock(clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_clock),
		.auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_reset(clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_reset),
		.auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_clock(clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_clock),
		.auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_reset(clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_reset),
		.auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_clock(clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_clock),
		.auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_reset(clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_reset),
		.auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_clock(clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_clock),
		.auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_reset(clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_reset)
	);
	ClockGroupResetSynchronizer resetSynchronizer(
		.auto_in_member_allClocks_implicit_clock_clock(resetSynchronizer_auto_in_member_allClocks_implicit_clock_clock),
		.auto_in_member_allClocks_implicit_clock_reset(resetSynchronizer_auto_in_member_allClocks_implicit_clock_reset),
		.auto_in_member_allClocks_subsystem_cbus_0_clock(resetSynchronizer_auto_in_member_allClocks_subsystem_cbus_0_clock),
		.auto_in_member_allClocks_subsystem_cbus_0_reset(resetSynchronizer_auto_in_member_allClocks_subsystem_cbus_0_reset),
		.auto_in_member_allClocks_subsystem_fbus_0_clock(resetSynchronizer_auto_in_member_allClocks_subsystem_fbus_0_clock),
		.auto_in_member_allClocks_subsystem_fbus_0_reset(resetSynchronizer_auto_in_member_allClocks_subsystem_fbus_0_reset),
		.auto_in_member_allClocks_subsystem_pbus_0_clock(resetSynchronizer_auto_in_member_allClocks_subsystem_pbus_0_clock),
		.auto_in_member_allClocks_subsystem_pbus_0_reset(resetSynchronizer_auto_in_member_allClocks_subsystem_pbus_0_reset),
		.auto_in_member_allClocks_subsystem_sbus_0_clock(resetSynchronizer_auto_in_member_allClocks_subsystem_sbus_0_clock),
		.auto_in_member_allClocks_subsystem_sbus_0_reset(resetSynchronizer_auto_in_member_allClocks_subsystem_sbus_0_reset),
		.auto_out_member_allClocks_implicit_clock_clock(resetSynchronizer_auto_out_member_allClocks_implicit_clock_clock),
		.auto_out_member_allClocks_implicit_clock_reset(resetSynchronizer_auto_out_member_allClocks_implicit_clock_reset),
		.auto_out_member_allClocks_subsystem_cbus_0_clock(resetSynchronizer_auto_out_member_allClocks_subsystem_cbus_0_clock),
		.auto_out_member_allClocks_subsystem_cbus_0_reset(resetSynchronizer_auto_out_member_allClocks_subsystem_cbus_0_reset),
		.auto_out_member_allClocks_subsystem_fbus_0_clock(resetSynchronizer_auto_out_member_allClocks_subsystem_fbus_0_clock),
		.auto_out_member_allClocks_subsystem_fbus_0_reset(resetSynchronizer_auto_out_member_allClocks_subsystem_fbus_0_reset),
		.auto_out_member_allClocks_subsystem_pbus_0_clock(resetSynchronizer_auto_out_member_allClocks_subsystem_pbus_0_clock),
		.auto_out_member_allClocks_subsystem_pbus_0_reset(resetSynchronizer_auto_out_member_allClocks_subsystem_pbus_0_reset),
		.auto_out_member_allClocks_subsystem_sbus_0_clock(resetSynchronizer_auto_out_member_allClocks_subsystem_sbus_0_clock),
		.auto_out_member_allClocks_subsystem_sbus_0_reset(resetSynchronizer_auto_out_member_allClocks_subsystem_sbus_0_reset)
	);
	ClockGroup_4 implicitClockGrouper(
		.auto_in_member_implicitClockGrouper_implicit_clock_clock(implicitClockGrouper_auto_in_member_implicitClockGrouper_implicit_clock_clock),
		.auto_in_member_implicitClockGrouper_implicit_clock_reset(implicitClockGrouper_auto_in_member_implicitClockGrouper_implicit_clock_reset),
		.auto_out_clock(implicitClockGrouper_auto_out_clock),
		.auto_out_reset(implicitClockGrouper_auto_out_reset)
	);
	DebugTransportModuleJTAG dtm(
		.io_jtag_clock(dtm_io_jtag_clock),
		.io_jtag_reset(dtm_io_jtag_reset),
		.io_dmi_req_ready(dtm_io_dmi_req_ready),
		.io_dmi_req_valid(dtm_io_dmi_req_valid),
		.io_dmi_req_bits_addr(dtm_io_dmi_req_bits_addr),
		.io_dmi_req_bits_data(dtm_io_dmi_req_bits_data),
		.io_dmi_req_bits_op(dtm_io_dmi_req_bits_op),
		.io_dmi_resp_ready(dtm_io_dmi_resp_ready),
		.io_dmi_resp_valid(dtm_io_dmi_resp_valid),
		.io_dmi_resp_bits_data(dtm_io_dmi_resp_bits_data),
		.io_dmi_resp_bits_resp(dtm_io_dmi_resp_bits_resp),
		.io_jtag_TMS(dtm_io_jtag_TMS),
		.io_jtag_TDI(dtm_io_jtag_TDI),
		.io_jtag_TDO_data(dtm_io_jtag_TDO_data)
	);
	assign auto_implicitClockGrouper_out_clock = implicitClockGrouper_auto_out_clock;
	assign auto_implicitClockGrouper_out_reset = implicitClockGrouper_auto_out_reset;
	assign auto_subsystem_cbus_fixedClockNode_out_clock = subsystem_cbus_auto_fixedClockNode_out_4_clock;
	assign auto_subsystem_cbus_fixedClockNode_out_reset = subsystem_cbus_auto_fixedClockNode_out_4_reset;
	assign serial_tl_clock = domain_clock;
	assign serial_tl_bits_in_ready = domain_serial_tl_in_ready;
	assign serial_tl_bits_out_valid = domain_serial_tl_out_valid;
	assign serial_tl_bits_out_bits = domain_serial_tl_out_bits;
	assign debug_systemjtag_jtag_TDO_data = dtm_io_jtag_TDO_data;
	assign debug_dmactive = debug_1_io_ctrl_dmactive;
	assign uart_0_txd = uartClockDomainWrapper_auto_uart_0_io_out_txd;
	assign ibus_auto_int_bus_int_in_0 = intsink_4_auto_out_0;
	assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_valid = tile_prci_domain_auto_tl_master_clock_xing_out_a_valid;
	assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode = tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_opcode;
	assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param = tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_param;
	assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size = tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_size;
	assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source = tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_source;
	assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address = tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_address;
	assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask = tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_mask;
	assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data = tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_data;
	assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_corrupt = tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_corrupt;
	assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_ready = tile_prci_domain_auto_tl_master_clock_xing_out_d_ready;
	assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid = subsystem_fbus_auto_bus_xing_out_a_valid;
	assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode = subsystem_fbus_auto_bus_xing_out_a_bits_opcode;
	assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param = subsystem_fbus_auto_bus_xing_out_a_bits_param;
	assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size = subsystem_fbus_auto_bus_xing_out_a_bits_size;
	assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source = subsystem_fbus_auto_bus_xing_out_a_bits_source;
	assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address = subsystem_fbus_auto_bus_xing_out_a_bits_address;
	assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask = subsystem_fbus_auto_bus_xing_out_a_bits_mask;
	assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data = subsystem_fbus_auto_bus_xing_out_a_bits_data;
	assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_corrupt = subsystem_fbus_auto_bus_xing_out_a_bits_corrupt;
	assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready = subsystem_fbus_auto_bus_xing_out_d_ready;
	assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready = subsystem_cbus_auto_bus_xing_in_a_ready;
	assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid = subsystem_cbus_auto_bus_xing_in_d_valid;
	assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode = subsystem_cbus_auto_bus_xing_in_d_bits_opcode;
	assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param = subsystem_cbus_auto_bus_xing_in_d_bits_param;
	assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size = subsystem_cbus_auto_bus_xing_in_d_bits_size;
	assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source = subsystem_cbus_auto_bus_xing_in_d_bits_source;
	assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink = subsystem_cbus_auto_bus_xing_in_d_bits_sink;
	assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied = subsystem_cbus_auto_bus_xing_in_d_bits_denied;
	assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data = subsystem_cbus_auto_bus_xing_in_d_bits_data;
	assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt = subsystem_cbus_auto_bus_xing_in_d_bits_corrupt;
	assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock = clockNamePrefixer_auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_clock;
	assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset = clockNamePrefixer_auto_clock_name_prefixer_out_0_member_subsystem_sbus_0_reset;
	assign subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_ready = uartClockDomainWrapper_auto_uart_0_control_xing_in_a_ready;
	assign subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_valid = uartClockDomainWrapper_auto_uart_0_control_xing_in_d_valid;
	assign subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode = uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_opcode;
	assign subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size = uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_size;
	assign subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source = uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_source;
	assign subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data = uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_data;
	assign subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_ready = domain_auto_tlserial_manager_crossing_in_a_ready;
	assign subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_valid = domain_auto_tlserial_manager_crossing_in_d_valid;
	assign subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_opcode = domain_auto_tlserial_manager_crossing_in_d_bits_opcode;
	assign subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_param = domain_auto_tlserial_manager_crossing_in_d_bits_param;
	assign subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_size = domain_auto_tlserial_manager_crossing_in_d_bits_size;
	assign subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_source = domain_auto_tlserial_manager_crossing_in_d_bits_source;
	assign subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_sink = domain_auto_tlserial_manager_crossing_in_d_bits_sink;
	assign subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_denied = domain_auto_tlserial_manager_crossing_in_d_bits_denied;
	assign subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_data = domain_auto_tlserial_manager_crossing_in_d_bits_data;
	assign subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_bits_corrupt = domain_auto_tlserial_manager_crossing_in_d_bits_corrupt;
	assign subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock = clockNamePrefixer_auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_clock;
	assign subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset = clockNamePrefixer_auto_clock_name_prefixer_out_1_member_subsystem_pbus_0_reset;
	assign subsystem_pbus_auto_bus_xing_in_a_valid = subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid;
	assign subsystem_pbus_auto_bus_xing_in_a_bits_opcode = subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode;
	assign subsystem_pbus_auto_bus_xing_in_a_bits_param = subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param;
	assign subsystem_pbus_auto_bus_xing_in_a_bits_size = subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size;
	assign subsystem_pbus_auto_bus_xing_in_a_bits_source = subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source;
	assign subsystem_pbus_auto_bus_xing_in_a_bits_address = subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address;
	assign subsystem_pbus_auto_bus_xing_in_a_bits_mask = subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask;
	assign subsystem_pbus_auto_bus_xing_in_a_bits_data = subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data;
	assign subsystem_pbus_auto_bus_xing_in_a_bits_corrupt = subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_corrupt;
	assign subsystem_pbus_auto_bus_xing_in_d_ready = subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready;
	assign subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_valid = domain_auto_serdesser_client_out_a_valid;
	assign subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_opcode = domain_auto_serdesser_client_out_a_bits_opcode;
	assign subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_param = domain_auto_serdesser_client_out_a_bits_param;
	assign subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_size = domain_auto_serdesser_client_out_a_bits_size;
	assign subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_source = domain_auto_serdesser_client_out_a_bits_source;
	assign subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_address = domain_auto_serdesser_client_out_a_bits_address;
	assign subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_mask = domain_auto_serdesser_client_out_a_bits_mask;
	assign subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_data = domain_auto_serdesser_client_out_a_bits_data;
	assign subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_bits_corrupt = domain_auto_serdesser_client_out_a_bits_corrupt;
	assign subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_ready = domain_auto_serdesser_client_out_d_ready;
	assign subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock = clockNamePrefixer_auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_clock;
	assign subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset = clockNamePrefixer_auto_clock_name_prefixer_out_2_member_subsystem_fbus_0_reset;
	assign subsystem_fbus_auto_bus_xing_out_a_ready = subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready;
	assign subsystem_fbus_auto_bus_xing_out_d_valid = subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid;
	assign subsystem_fbus_auto_bus_xing_out_d_bits_opcode = subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode;
	assign subsystem_fbus_auto_bus_xing_out_d_bits_param = subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param;
	assign subsystem_fbus_auto_bus_xing_out_d_bits_size = subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size;
	assign subsystem_fbus_auto_bus_xing_out_d_bits_sink = subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink;
	assign subsystem_fbus_auto_bus_xing_out_d_bits_denied = subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied;
	assign subsystem_fbus_auto_bus_xing_out_d_bits_data = subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data;
	assign subsystem_fbus_auto_bus_xing_out_d_bits_corrupt = subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt;
	assign subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_ready = prci_ctrl_domain_auto_tileResetSetter_tl_in_a_ready;
	assign subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_valid = prci_ctrl_domain_auto_tileResetSetter_tl_in_d_valid;
	assign subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_opcode = prci_ctrl_domain_auto_tileResetSetter_tl_in_d_bits_opcode;
	assign subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_size = prci_ctrl_domain_auto_tileResetSetter_tl_in_d_bits_size;
	assign subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_source = prci_ctrl_domain_auto_tileResetSetter_tl_in_d_bits_source;
	assign subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_bits_data = prci_ctrl_domain_auto_tileResetSetter_tl_in_d_bits_data;
	assign subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_ready = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_ready;
	assign subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_valid = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_valid;
	assign subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_opcode = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_bits_opcode;
	assign subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_size = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_bits_size;
	assign subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_source = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_bits_source;
	assign subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_bits_data = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_bits_data;
	assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_ready = bootROMDomainWrapper_auto_bootrom_in_a_ready;
	assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_valid = bootROMDomainWrapper_auto_bootrom_in_d_valid;
	assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_size = bootROMDomainWrapper_auto_bootrom_in_d_bits_size;
	assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_source = bootROMDomainWrapper_auto_bootrom_in_d_bits_source;
	assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_data = bootROMDomainWrapper_auto_bootrom_in_d_bits_data;
	assign subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_ready = tile_prci_domain_auto_tl_slave_clock_xing_in_a_ready;
	assign subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_valid = tile_prci_domain_auto_tl_slave_clock_xing_in_d_valid;
	assign subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_opcode = tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_opcode;
	assign subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_param = tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_param;
	assign subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_size = tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_size;
	assign subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_source = tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_source;
	assign subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_sink = tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_sink;
	assign subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_denied = tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_denied;
	assign subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_data = tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_data;
	assign subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_bits_corrupt = tile_prci_domain_auto_tl_slave_clock_xing_in_d_bits_corrupt;
	assign subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_ready = debug_1_auto_dmInner_dmInner_tl_in_a_ready;
	assign subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_valid = debug_1_auto_dmInner_dmInner_tl_in_d_valid;
	assign subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_bits_opcode = debug_1_auto_dmInner_dmInner_tl_in_d_bits_opcode;
	assign subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_bits_size = debug_1_auto_dmInner_dmInner_tl_in_d_bits_size;
	assign subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_bits_source = debug_1_auto_dmInner_dmInner_tl_in_d_bits_source;
	assign subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_bits_data = debug_1_auto_dmInner_dmInner_tl_in_d_bits_data;
	assign subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_ready = clint_auto_in_a_ready;
	assign subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_valid = clint_auto_in_d_valid;
	assign subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_opcode = clint_auto_in_d_bits_opcode;
	assign subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_size = clint_auto_in_d_bits_size;
	assign subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_source = clint_auto_in_d_bits_source;
	assign subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_data = clint_auto_in_d_bits_data;
	assign subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_ready = plicDomainWrapper_auto_plic_in_a_ready;
	assign subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_valid = plicDomainWrapper_auto_plic_in_d_valid;
	assign subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_opcode = plicDomainWrapper_auto_plic_in_d_bits_opcode;
	assign subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_size = plicDomainWrapper_auto_plic_in_d_bits_size;
	assign subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_source = plicDomainWrapper_auto_plic_in_d_bits_source;
	assign subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_data = plicDomainWrapper_auto_plic_in_d_bits_data;
	assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready = subsystem_pbus_auto_bus_xing_in_a_ready;
	assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid = subsystem_pbus_auto_bus_xing_in_d_valid;
	assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode = subsystem_pbus_auto_bus_xing_in_d_bits_opcode;
	assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_param = subsystem_pbus_auto_bus_xing_in_d_bits_param;
	assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size = subsystem_pbus_auto_bus_xing_in_d_bits_size;
	assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source = subsystem_pbus_auto_bus_xing_in_d_bits_source;
	assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_sink = subsystem_pbus_auto_bus_xing_in_d_bits_sink;
	assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied = subsystem_pbus_auto_bus_xing_in_d_bits_denied;
	assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data = subsystem_pbus_auto_bus_xing_in_d_bits_data;
	assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt = subsystem_pbus_auto_bus_xing_in_d_bits_corrupt;
	assign subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock = clockNamePrefixer_auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_clock;
	assign subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset = clockNamePrefixer_auto_clock_name_prefixer_out_3_member_subsystem_cbus_0_reset;
	assign subsystem_cbus_auto_bus_xing_in_a_valid = subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid;
	assign subsystem_cbus_auto_bus_xing_in_a_bits_opcode = subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode;
	assign subsystem_cbus_auto_bus_xing_in_a_bits_param = subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param;
	assign subsystem_cbus_auto_bus_xing_in_a_bits_size = subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size;
	assign subsystem_cbus_auto_bus_xing_in_a_bits_source = subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source;
	assign subsystem_cbus_auto_bus_xing_in_a_bits_address = subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address;
	assign subsystem_cbus_auto_bus_xing_in_a_bits_mask = subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask;
	assign subsystem_cbus_auto_bus_xing_in_a_bits_data = subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data;
	assign subsystem_cbus_auto_bus_xing_in_a_bits_corrupt = subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt;
	assign subsystem_cbus_auto_bus_xing_in_d_ready = subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready;
	assign subsystem_cbus_custom_boot = custom_boot;
	assign tile_prci_domain_auto_intsink_in_sync_0 = debug_1_auto_dmOuter_intsource_out_sync_0;
	assign tile_prci_domain_auto_tile_reset_domain_tile_hartid_in = tileHartIdNexusNode_auto_out;
	assign tile_prci_domain_auto_int_in_clock_xing_in_1_sync_0 = intsource_1_auto_out_sync_0;
	assign tile_prci_domain_auto_int_in_clock_xing_in_0_sync_0 = intsource_auto_out_sync_0;
	assign tile_prci_domain_auto_int_in_clock_xing_in_0_sync_1 = intsource_auto_out_sync_1;
	assign tile_prci_domain_auto_tl_slave_clock_xing_in_a_valid = subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_valid;
	assign tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_opcode = subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_opcode;
	assign tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_param = subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_param;
	assign tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_size = subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_size;
	assign tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_source = subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_source;
	assign tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_address = subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_address;
	assign tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_mask = subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_mask;
	assign tile_prci_domain_auto_tl_slave_clock_xing_in_a_bits_data = subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_a_bits_data;
	assign tile_prci_domain_auto_tl_slave_clock_xing_in_d_ready = subsystem_cbus_auto_coupler_to_tile_tl_slave_clock_xing_out_d_ready;
	assign tile_prci_domain_auto_tl_master_clock_xing_out_a_ready = subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_ready;
	assign tile_prci_domain_auto_tl_master_clock_xing_out_d_valid = subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_valid;
	assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_opcode = subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode;
	assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_param = subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param;
	assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_size = subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size;
	assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_source = subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source;
	assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_sink = subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink;
	assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_denied = subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied;
	assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_data = subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data;
	assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_corrupt = subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt;
	assign tile_prci_domain_auto_tap_clock_in_clock = subsystem_sbus_auto_fixedClockNode_out_1_clock;
	assign tile_prci_domain_auto_tap_clock_in_reset = subsystem_sbus_auto_fixedClockNode_out_1_reset;
	assign plicDomainWrapper_auto_plic_int_in_0 = ibus_auto_int_bus_int_out_0;
	assign plicDomainWrapper_auto_plic_in_a_valid = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_valid;
	assign plicDomainWrapper_auto_plic_in_a_bits_opcode = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_opcode;
	assign plicDomainWrapper_auto_plic_in_a_bits_param = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_param;
	assign plicDomainWrapper_auto_plic_in_a_bits_size = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_size;
	assign plicDomainWrapper_auto_plic_in_a_bits_source = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_source;
	assign plicDomainWrapper_auto_plic_in_a_bits_address = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_address;
	assign plicDomainWrapper_auto_plic_in_a_bits_mask = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_mask;
	assign plicDomainWrapper_auto_plic_in_a_bits_data = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_data;
	assign plicDomainWrapper_auto_plic_in_a_bits_corrupt = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_corrupt;
	assign plicDomainWrapper_auto_plic_in_d_ready = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_ready;
	assign plicDomainWrapper_auto_clock_in_clock = subsystem_cbus_auto_fixedClockNode_out_0_clock;
	assign plicDomainWrapper_auto_clock_in_reset = subsystem_cbus_auto_fixedClockNode_out_0_reset;
	assign clint_clock = subsystem_cbus_clock;
	assign clint_reset = subsystem_cbus_reset;
	assign clint_auto_in_a_valid = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_valid;
	assign clint_auto_in_a_bits_opcode = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_opcode;
	assign clint_auto_in_a_bits_param = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_param;
	assign clint_auto_in_a_bits_size = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_size;
	assign clint_auto_in_a_bits_source = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_source;
	assign clint_auto_in_a_bits_address = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_address;
	assign clint_auto_in_a_bits_mask = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_mask;
	assign clint_auto_in_a_bits_data = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_data;
	assign clint_auto_in_a_bits_corrupt = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_corrupt;
	assign clint_auto_in_d_ready = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_ready;
	assign clint_io_rtcTick = int_rtc_tick_value == 7'h63;
	assign debug_1_auto_dmInner_dmInner_tl_in_a_valid = subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_valid;
	assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_opcode = subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_opcode;
	assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_param = subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_param;
	assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_size = subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_size;
	assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_source = subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_source;
	assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_address = subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_address;
	assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_mask = subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_mask;
	assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_data = subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_data;
	assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_corrupt = subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_corrupt;
	assign debug_1_auto_dmInner_dmInner_tl_in_d_ready = subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_ready;
	assign debug_1_io_debug_clock = debug_clock;
	assign debug_1_io_debug_reset = debug_reset;
	assign debug_1_io_ctrl_dmactiveAck = debug_dmactiveAck;
	assign debug_1_io_dmi_dmi_req_valid = dtm_io_dmi_req_valid;
	assign debug_1_io_dmi_dmi_req_bits_addr = dtm_io_dmi_req_bits_addr;
	assign debug_1_io_dmi_dmi_req_bits_data = dtm_io_dmi_req_bits_data;
	assign debug_1_io_dmi_dmi_req_bits_op = dtm_io_dmi_req_bits_op;
	assign debug_1_io_dmi_dmi_resp_ready = dtm_io_dmi_resp_ready;
	assign debug_1_io_dmi_dmiClock = debug_systemjtag_jtag_TCK;
	assign debug_1_io_dmi_dmiReset = debug_systemjtag_reset;
	assign debug_1_io_hartIsInReset_0 = resetctrl_hartIsInReset_0;
	assign xbar_auto_int_in_0 = intsink_1_auto_out_0;
	assign xbar_1_auto_int_in_0 = intsink_2_auto_out_0;
	assign xbar_2_auto_int_in_0 = intsink_3_auto_out_0;
	assign intsource_clock = clock;
	assign intsource_reset = reset;
	assign intsource_auto_in_0 = clint_auto_int_out_0;
	assign intsource_auto_in_1 = clint_auto_int_out_1;
	assign intsource_1_clock = clock;
	assign intsource_1_reset = reset;
	assign intsource_1_auto_in_0 = plicDomainWrapper_auto_plic_int_out_0;
	assign intsink_1_auto_in_sync_0 = tile_prci_domain_auto_int_out_clock_xing_out_0_sync_0;
	assign intsink_2_auto_in_sync_0 = tile_prci_domain_auto_int_out_clock_xing_out_1_sync_0;
	assign intsink_3_auto_in_sync_0 = tile_prci_domain_auto_int_out_clock_xing_out_2_sync_0;
	assign bootROMDomainWrapper_auto_bootrom_in_a_valid = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_valid;
	assign bootROMDomainWrapper_auto_bootrom_in_a_bits_opcode = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode;
	assign bootROMDomainWrapper_auto_bootrom_in_a_bits_param = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_param;
	assign bootROMDomainWrapper_auto_bootrom_in_a_bits_size = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_size;
	assign bootROMDomainWrapper_auto_bootrom_in_a_bits_source = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_source;
	assign bootROMDomainWrapper_auto_bootrom_in_a_bits_address = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_address;
	assign bootROMDomainWrapper_auto_bootrom_in_a_bits_mask = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_mask;
	assign bootROMDomainWrapper_auto_bootrom_in_a_bits_corrupt = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt;
	assign bootROMDomainWrapper_auto_bootrom_in_d_ready = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_ready;
	assign bootROMDomainWrapper_auto_clock_in_clock = subsystem_cbus_auto_fixedClockNode_out_2_clock;
	assign bootROMDomainWrapper_auto_clock_in_reset = subsystem_cbus_auto_fixedClockNode_out_2_reset;
	assign domain_auto_serdesser_client_out_a_ready = subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_a_ready;
	assign domain_auto_serdesser_client_out_d_valid = subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_valid;
	assign domain_auto_serdesser_client_out_d_bits_opcode = subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_opcode;
	assign domain_auto_serdesser_client_out_d_bits_param = subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_param;
	assign domain_auto_serdesser_client_out_d_bits_size = subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_size;
	assign domain_auto_serdesser_client_out_d_bits_source = subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_source;
	assign domain_auto_serdesser_client_out_d_bits_sink = subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_sink;
	assign domain_auto_serdesser_client_out_d_bits_denied = subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_denied;
	assign domain_auto_serdesser_client_out_d_bits_data = subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_data;
	assign domain_auto_serdesser_client_out_d_bits_corrupt = subsystem_fbus_auto_coupler_from_port_named_serial_tl_ctrl_buffer_in_d_bits_corrupt;
	assign domain_auto_tlserial_manager_crossing_in_a_valid = subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_valid;
	assign domain_auto_tlserial_manager_crossing_in_a_bits_opcode = subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_opcode;
	assign domain_auto_tlserial_manager_crossing_in_a_bits_param = subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_param;
	assign domain_auto_tlserial_manager_crossing_in_a_bits_size = subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_size;
	assign domain_auto_tlserial_manager_crossing_in_a_bits_source = subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_source;
	assign domain_auto_tlserial_manager_crossing_in_a_bits_address = subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_address;
	assign domain_auto_tlserial_manager_crossing_in_a_bits_mask = subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_mask;
	assign domain_auto_tlserial_manager_crossing_in_a_bits_data = subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_data;
	assign domain_auto_tlserial_manager_crossing_in_a_bits_corrupt = subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_a_bits_corrupt;
	assign domain_auto_tlserial_manager_crossing_in_d_ready = subsystem_pbus_auto_coupler_to_port_named_serial_tl_mem_tlserial_manager_crossing_out_d_ready;
	assign domain_auto_clock_in_clock = subsystem_fbus_auto_fixedClockNode_out_clock;
	assign domain_auto_clock_in_reset = subsystem_fbus_auto_fixedClockNode_out_reset;
	assign domain_serial_tl_in_valid = serial_tl_bits_in_valid;
	assign domain_serial_tl_in_bits = serial_tl_bits_in_bits;
	assign domain_serial_tl_out_ready = serial_tl_bits_out_ready;
	assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_valid = subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_valid;
	assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_opcode = subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode;
	assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_param = subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_param;
	assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_size = subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size;
	assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_source = subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source;
	assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_address = subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address;
	assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_mask = subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask;
	assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_data = subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data;
	assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_corrupt = subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_corrupt;
	assign uartClockDomainWrapper_auto_uart_0_control_xing_in_d_ready = subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_ready;
	assign uartClockDomainWrapper_auto_uart_0_io_out_rxd = uart_0_rxd;
	assign uartClockDomainWrapper_auto_clock_in_clock = subsystem_pbus_auto_fixedClockNode_out_clock;
	assign uartClockDomainWrapper_auto_clock_in_reset = subsystem_pbus_auto_fixedClockNode_out_reset;
	assign intsink_4_auto_in_sync_0 = uartClockDomainWrapper_auto_uart_0_int_xing_out_sync_0;
	assign prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock = auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock;
	assign prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset = auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset;
	assign prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock = auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock;
	assign prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset = auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset;
	assign prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock = auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock;
	assign prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset = auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset;
	assign prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock = auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock;
	assign prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset = auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset;
	assign prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock = auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock;
	assign prci_ctrl_domain_auto_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset = auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset;
	assign prci_ctrl_domain_auto_tileResetSetter_tl_in_a_valid = subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_valid;
	assign prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_opcode = subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_opcode;
	assign prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_param = subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_param;
	assign prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_size = subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_size;
	assign prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_source = subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_source;
	assign prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_address = subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_address;
	assign prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_mask = subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_mask;
	assign prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_data = subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_data;
	assign prci_ctrl_domain_auto_tileResetSetter_tl_in_a_bits_corrupt = subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_a_bits_corrupt;
	assign prci_ctrl_domain_auto_tileResetSetter_tl_in_d_ready = subsystem_cbus_auto_coupler_to_slave_named_tileresetsetter_buffer_out_d_ready;
	assign prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_valid = subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_valid;
	assign prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_opcode = subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_opcode;
	assign prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_param = subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_param;
	assign prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_size = subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_size;
	assign prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_source = subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_source;
	assign prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_address = subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_address;
	assign prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_mask = subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_mask;
	assign prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_data = subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_data;
	assign prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_a_bits_corrupt = subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_a_bits_corrupt;
	assign prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_in_d_ready = subsystem_cbus_auto_coupler_to_slave_named_clockgater_buffer_out_d_ready;
	assign prci_ctrl_domain_auto_clock_in_clock = subsystem_cbus_auto_fixedClockNode_out_3_clock;
	assign prci_ctrl_domain_auto_clock_in_reset = subsystem_cbus_auto_fixedClockNode_out_3_reset;
	assign aggregator_auto_in_member_allClocks_implicit_clock_clock = frequencySpecifier_auto_frequency_specifier_out_member_allClocks_implicit_clock_clock;
	assign aggregator_auto_in_member_allClocks_implicit_clock_reset = frequencySpecifier_auto_frequency_specifier_out_member_allClocks_implicit_clock_reset;
	assign aggregator_auto_in_member_allClocks_subsystem_cbus_0_clock = frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_clock;
	assign aggregator_auto_in_member_allClocks_subsystem_cbus_0_reset = frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_cbus_0_reset;
	assign aggregator_auto_in_member_allClocks_subsystem_fbus_0_clock = frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_clock;
	assign aggregator_auto_in_member_allClocks_subsystem_fbus_0_reset = frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_fbus_0_reset;
	assign aggregator_auto_in_member_allClocks_subsystem_pbus_0_clock = frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_clock;
	assign aggregator_auto_in_member_allClocks_subsystem_pbus_0_reset = frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_pbus_0_reset;
	assign aggregator_auto_in_member_allClocks_subsystem_sbus_0_clock = frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_clock;
	assign aggregator_auto_in_member_allClocks_subsystem_sbus_0_reset = frequencySpecifier_auto_frequency_specifier_out_member_allClocks_subsystem_sbus_0_reset;
	assign clockNamePrefixer_auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_clock = aggregator_auto_out_3_member_subsystem_cbus_subsystem_cbus_0_clock;
	assign clockNamePrefixer_auto_clock_name_prefixer_in_3_member_subsystem_cbus_subsystem_cbus_0_reset = aggregator_auto_out_3_member_subsystem_cbus_subsystem_cbus_0_reset;
	assign clockNamePrefixer_auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_clock = aggregator_auto_out_2_member_subsystem_fbus_subsystem_fbus_0_clock;
	assign clockNamePrefixer_auto_clock_name_prefixer_in_2_member_subsystem_fbus_subsystem_fbus_0_reset = aggregator_auto_out_2_member_subsystem_fbus_subsystem_fbus_0_reset;
	assign clockNamePrefixer_auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_clock = aggregator_auto_out_1_member_subsystem_pbus_subsystem_pbus_0_clock;
	assign clockNamePrefixer_auto_clock_name_prefixer_in_1_member_subsystem_pbus_subsystem_pbus_0_reset = aggregator_auto_out_1_member_subsystem_pbus_subsystem_pbus_0_reset;
	assign clockNamePrefixer_auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_clock = aggregator_auto_out_0_member_subsystem_sbus_subsystem_sbus_0_clock;
	assign clockNamePrefixer_auto_clock_name_prefixer_in_0_member_subsystem_sbus_subsystem_sbus_0_reset = aggregator_auto_out_0_member_subsystem_sbus_subsystem_sbus_0_reset;
	assign frequencySpecifier_auto_frequency_specifier_in_member_allClocks_implicit_clock_clock = clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_implicit_clock_clock;
	assign frequencySpecifier_auto_frequency_specifier_in_member_allClocks_implicit_clock_reset = clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_implicit_clock_reset;
	assign frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_clock = clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_clock;
	assign frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_cbus_0_reset = clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_cbus_0_reset;
	assign frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_clock = clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_clock;
	assign frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_fbus_0_reset = clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_fbus_0_reset;
	assign frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_clock = clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_clock;
	assign frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_pbus_0_reset = clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_pbus_0_reset;
	assign frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_clock = clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_clock;
	assign frequencySpecifier_auto_frequency_specifier_in_member_allClocks_subsystem_sbus_0_reset = clockGroupCombiner_auto_clock_group_combiner_out_member_allClocks_subsystem_sbus_0_reset;
	assign clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_implicit_clock_clock = resetSynchronizer_auto_out_member_allClocks_implicit_clock_clock;
	assign clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_implicit_clock_reset = resetSynchronizer_auto_out_member_allClocks_implicit_clock_reset;
	assign clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_clock = resetSynchronizer_auto_out_member_allClocks_subsystem_cbus_0_clock;
	assign clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_cbus_0_reset = resetSynchronizer_auto_out_member_allClocks_subsystem_cbus_0_reset;
	assign clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_clock = resetSynchronizer_auto_out_member_allClocks_subsystem_fbus_0_clock;
	assign clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_fbus_0_reset = resetSynchronizer_auto_out_member_allClocks_subsystem_fbus_0_reset;
	assign clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_clock = resetSynchronizer_auto_out_member_allClocks_subsystem_pbus_0_clock;
	assign clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_pbus_0_reset = resetSynchronizer_auto_out_member_allClocks_subsystem_pbus_0_reset;
	assign clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_clock = resetSynchronizer_auto_out_member_allClocks_subsystem_sbus_0_clock;
	assign clockGroupCombiner_auto_clock_group_combiner_in_member_allClocks_subsystem_sbus_0_reset = resetSynchronizer_auto_out_member_allClocks_subsystem_sbus_0_reset;
	assign resetSynchronizer_auto_in_member_allClocks_implicit_clock_clock = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_clock;
	assign resetSynchronizer_auto_in_member_allClocks_implicit_clock_reset = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_implicit_clock_reset;
	assign resetSynchronizer_auto_in_member_allClocks_subsystem_cbus_0_clock = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_clock;
	assign resetSynchronizer_auto_in_member_allClocks_subsystem_cbus_0_reset = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_cbus_0_reset;
	assign resetSynchronizer_auto_in_member_allClocks_subsystem_fbus_0_clock = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_clock;
	assign resetSynchronizer_auto_in_member_allClocks_subsystem_fbus_0_reset = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_fbus_0_reset;
	assign resetSynchronizer_auto_in_member_allClocks_subsystem_pbus_0_clock = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_clock;
	assign resetSynchronizer_auto_in_member_allClocks_subsystem_pbus_0_reset = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_pbus_0_reset;
	assign resetSynchronizer_auto_in_member_allClocks_subsystem_sbus_0_clock = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_clock;
	assign resetSynchronizer_auto_in_member_allClocks_subsystem_sbus_0_reset = prci_ctrl_domain_auto_tileClockGater_tile_clock_gater_out_member_allClocks_subsystem_sbus_0_reset;
	assign implicitClockGrouper_auto_in_member_implicitClockGrouper_implicit_clock_clock = aggregator_auto_out_4_member_implicitClockGrouper_implicit_clock_clock;
	assign implicitClockGrouper_auto_in_member_implicitClockGrouper_implicit_clock_reset = aggregator_auto_out_4_member_implicitClockGrouper_implicit_clock_reset;
	assign dtm_io_jtag_clock = debug_systemjtag_jtag_TCK;
	assign dtm_io_jtag_reset = debug_systemjtag_reset;
	assign dtm_io_dmi_req_ready = debug_1_io_dmi_dmi_req_ready;
	assign dtm_io_dmi_resp_valid = debug_1_io_dmi_dmi_resp_valid;
	assign dtm_io_dmi_resp_bits_data = debug_1_io_dmi_dmi_resp_bits_data;
	assign dtm_io_dmi_resp_bits_resp = debug_1_io_dmi_dmi_resp_bits_resp;
	assign dtm_io_jtag_TMS = debug_systemjtag_jtag_TMS;
	assign dtm_io_jtag_TDI = debug_systemjtag_jtag_TDI;
	always @(posedge subsystem_pbus_clock)
		if (subsystem_pbus_reset)
			int_rtc_tick_value <= 7'h00;
		else if (int_rtc_tick_wrap_wrap)
			int_rtc_tick_value <= 7'h00;
		else
			int_rtc_tick_value <= _int_rtc_tick_wrap_value_T_1;
endmodule
module DividerOnlyClockGenerator (
	auto_divider_only_clock_gen_in_clock,
	auto_divider_only_clock_gen_in_reset,
	auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_clock,
	auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_reset,
	auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_clock,
	auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_reset,
	auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_clock,
	auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_reset,
	auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_clock,
	auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_reset,
	auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_clock,
	auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_reset
);
	input auto_divider_only_clock_gen_in_clock;
	input auto_divider_only_clock_gen_in_reset;
	output wire auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_clock;
	output wire auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_reset;
	output wire auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_clock;
	output wire auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_reset;
	output wire auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_clock;
	output wire auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_reset;
	output wire auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_clock;
	output wire auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_reset;
	output wire auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_clock;
	output wire auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_reset;
	wire bundleOut_0_member_allClocks_subsystem_sbus_0_clock_ClockDivideBy1_clk_out;
	wire bundleOut_0_member_allClocks_subsystem_sbus_0_clock_ClockDivideBy1_clk_in;
	ClockDividerN #(.DIV(1)) bundleOut_0_member_allClocks_subsystem_sbus_0_clock_ClockDivideBy1(
		.clk_out(bundleOut_0_member_allClocks_subsystem_sbus_0_clock_ClockDivideBy1_clk_out),
		.clk_in(bundleOut_0_member_allClocks_subsystem_sbus_0_clock_ClockDivideBy1_clk_in)
	);
	assign auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_clock = bundleOut_0_member_allClocks_subsystem_sbus_0_clock_ClockDivideBy1_clk_out;
	assign auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_reset = auto_divider_only_clock_gen_in_reset;
	assign auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_clock = bundleOut_0_member_allClocks_subsystem_sbus_0_clock_ClockDivideBy1_clk_out;
	assign auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_reset = auto_divider_only_clock_gen_in_reset;
	assign auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_clock = bundleOut_0_member_allClocks_subsystem_sbus_0_clock_ClockDivideBy1_clk_out;
	assign auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_reset = auto_divider_only_clock_gen_in_reset;
	assign auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_clock = bundleOut_0_member_allClocks_subsystem_sbus_0_clock_ClockDivideBy1_clk_out;
	assign auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_reset = auto_divider_only_clock_gen_in_reset;
	assign auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_clock = bundleOut_0_member_allClocks_subsystem_sbus_0_clock_ClockDivideBy1_clk_out;
	assign auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_reset = auto_divider_only_clock_gen_in_reset;
	assign bundleOut_0_member_allClocks_subsystem_sbus_0_clock_ClockDivideBy1_clk_in = auto_divider_only_clock_gen_in_clock;
endmodule
module ResetSynchronizerShiftReg_w1_d3_i0 (
	clock,
	reset,
	io_d,
	io_q
);
	input clock;
	input reset;
	input io_d;
	output wire io_q;
	wire output_chain_clock;
	wire output_chain_reset;
	wire output_chain_io_d;
	wire output_chain_io_q;
	AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain(
		.clock(output_chain_clock),
		.reset(output_chain_reset),
		.io_d(output_chain_io_d),
		.io_q(output_chain_io_q)
	);
	assign io_q = output_chain_io_q;
	assign output_chain_clock = clock;
	assign output_chain_reset = reset;
	assign output_chain_io_d = io_d;
endmodule
module ChipTop (
	vccd1,
	vssd1,
	jtag_TCK,
	jtag_TMS,
	jtag_TDI,
	jtag_TDO,
	serial_tl_clock,
	serial_tl_bits_in_ready,
	serial_tl_bits_in_valid,
	serial_tl_bits_in_bits,
	serial_tl_bits_out_ready,
	serial_tl_bits_out_valid,
	serial_tl_bits_out_bits,
	custom_boot,
	clock_clock,
	reset,
	uart_0_txd,
	uart_0_rxd
);
    inout vccd1;
	inout vssd1;
	input jtag_TCK;
	input jtag_TMS;
	input jtag_TDI;
	output wire jtag_TDO;
	output wire serial_tl_clock;
	output wire serial_tl_bits_in_ready;
	input serial_tl_bits_in_valid;
	input [31:0] serial_tl_bits_in_bits;
	input serial_tl_bits_out_ready;
	output wire serial_tl_bits_out_valid;
	output wire [31:0] serial_tl_bits_out_bits;
	input custom_boot;
	input clock_clock;
	input reset;
	output wire uart_0_txd;
	input uart_0_rxd;
	wire system_clock;
	wire system_reset;
	wire system_auto_implicitClockGrouper_out_clock;
	wire system_auto_implicitClockGrouper_out_reset;
	wire system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock;
	wire system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset;
	wire system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock;
	wire system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset;
	wire system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock;
	wire system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset;
	wire system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock;
	wire system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset;
	wire system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock;
	wire system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset;
	wire system_auto_subsystem_cbus_fixedClockNode_out_clock;
	wire system_auto_subsystem_cbus_fixedClockNode_out_reset;
	wire system_custom_boot;
	wire system_serial_tl_clock;
	wire system_serial_tl_bits_in_ready;
	wire system_serial_tl_bits_in_valid;
	wire [31:0] system_serial_tl_bits_in_bits;
	wire system_serial_tl_bits_out_ready;
	wire system_serial_tl_bits_out_valid;
	wire [31:0] system_serial_tl_bits_out_bits;
	wire system_resetctrl_hartIsInReset_0;
	wire system_debug_clock;
	wire system_debug_reset;
	wire system_debug_systemjtag_jtag_TCK;
	wire system_debug_systemjtag_jtag_TMS;
	wire system_debug_systemjtag_jtag_TDI;
	wire system_debug_systemjtag_jtag_TDO_data;
	wire system_debug_systemjtag_reset;
	wire system_debug_dmactive;
	wire system_debug_dmactiveAck;
	wire system_uart_0_txd;
	wire system_uart_0_rxd;
	wire dividerOnlyClockGen_auto_divider_only_clock_gen_in_clock;
	wire dividerOnlyClockGen_auto_divider_only_clock_gen_in_reset;
	wire dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_clock;
	wire dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_reset;
	wire dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_clock;
	wire dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_reset;
	wire dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_clock;
	wire dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_reset;
	wire dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_clock;
	wire dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_reset;
	wire dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_clock;
	wire dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_reset;
	wire system_debug_systemjtag_reset_catcher_clock;
	wire system_debug_systemjtag_reset_catcher_reset;
	wire system_debug_systemjtag_reset_catcher_io_sync_reset;
	wire debug_reset_syncd_debug_reset_sync_clock;
	wire debug_reset_syncd_debug_reset_sync_reset;
	wire debug_reset_syncd_debug_reset_sync_io_d;
	wire debug_reset_syncd_debug_reset_sync_io_q;
	wire dmactiveAck_dmactiveAck_clock;
	wire dmactiveAck_dmactiveAck_reset;
	wire dmactiveAck_dmactiveAck_io_d;
	wire dmactiveAck_dmactiveAck_io_q;
	wire gated_clock_debug_clock_gate_in;
	wire gated_clock_debug_clock_gate_test_en;
	wire gated_clock_debug_clock_gate_en;
	wire gated_clock_debug_clock_gate_out;
	wire iocell_jtag_TDO_pad;
	wire iocell_jtag_TDO_o;
	wire iocell_jtag_TDO_oe;
	wire iocell_jtag_TDI_pad;
	wire iocell_jtag_TDI_i;
	wire iocell_jtag_TDI_ie;
	wire iocell_jtag_TMS_pad;
	wire iocell_jtag_TMS_i;
	wire iocell_jtag_TMS_ie;
	wire iocell_jtag_TCK_pad;
	wire iocell_jtag_TCK_i;
	wire iocell_jtag_TCK_ie;
	wire iocell_serial_tl_bits_out_bits_pad;
	wire iocell_serial_tl_bits_out_bits_o;
	wire iocell_serial_tl_bits_out_bits_oe;
	wire iocell_serial_tl_bits_out_bits_1_pad;
	wire iocell_serial_tl_bits_out_bits_1_o;
	wire iocell_serial_tl_bits_out_bits_1_oe;
	wire iocell_serial_tl_bits_out_bits_2_pad;
	wire iocell_serial_tl_bits_out_bits_2_o;
	wire iocell_serial_tl_bits_out_bits_2_oe;
	wire iocell_serial_tl_bits_out_bits_3_pad;
	wire iocell_serial_tl_bits_out_bits_3_o;
	wire iocell_serial_tl_bits_out_bits_3_oe;
	wire iocell_serial_tl_bits_out_bits_4_pad;
	wire iocell_serial_tl_bits_out_bits_4_o;
	wire iocell_serial_tl_bits_out_bits_4_oe;
	wire iocell_serial_tl_bits_out_bits_5_pad;
	wire iocell_serial_tl_bits_out_bits_5_o;
	wire iocell_serial_tl_bits_out_bits_5_oe;
	wire iocell_serial_tl_bits_out_bits_6_pad;
	wire iocell_serial_tl_bits_out_bits_6_o;
	wire iocell_serial_tl_bits_out_bits_6_oe;
	wire iocell_serial_tl_bits_out_bits_7_pad;
	wire iocell_serial_tl_bits_out_bits_7_o;
	wire iocell_serial_tl_bits_out_bits_7_oe;
	wire iocell_serial_tl_bits_out_bits_8_pad;
	wire iocell_serial_tl_bits_out_bits_8_o;
	wire iocell_serial_tl_bits_out_bits_8_oe;
	wire iocell_serial_tl_bits_out_bits_9_pad;
	wire iocell_serial_tl_bits_out_bits_9_o;
	wire iocell_serial_tl_bits_out_bits_9_oe;
	wire iocell_serial_tl_bits_out_bits_10_pad;
	wire iocell_serial_tl_bits_out_bits_10_o;
	wire iocell_serial_tl_bits_out_bits_10_oe;
	wire iocell_serial_tl_bits_out_bits_11_pad;
	wire iocell_serial_tl_bits_out_bits_11_o;
	wire iocell_serial_tl_bits_out_bits_11_oe;
	wire iocell_serial_tl_bits_out_bits_12_pad;
	wire iocell_serial_tl_bits_out_bits_12_o;
	wire iocell_serial_tl_bits_out_bits_12_oe;
	wire iocell_serial_tl_bits_out_bits_13_pad;
	wire iocell_serial_tl_bits_out_bits_13_o;
	wire iocell_serial_tl_bits_out_bits_13_oe;
	wire iocell_serial_tl_bits_out_bits_14_pad;
	wire iocell_serial_tl_bits_out_bits_14_o;
	wire iocell_serial_tl_bits_out_bits_14_oe;
	wire iocell_serial_tl_bits_out_bits_15_pad;
	wire iocell_serial_tl_bits_out_bits_15_o;
	wire iocell_serial_tl_bits_out_bits_15_oe;
	wire iocell_serial_tl_bits_out_bits_16_pad;
	wire iocell_serial_tl_bits_out_bits_16_o;
	wire iocell_serial_tl_bits_out_bits_16_oe;
	wire iocell_serial_tl_bits_out_bits_17_pad;
	wire iocell_serial_tl_bits_out_bits_17_o;
	wire iocell_serial_tl_bits_out_bits_17_oe;
	wire iocell_serial_tl_bits_out_bits_18_pad;
	wire iocell_serial_tl_bits_out_bits_18_o;
	wire iocell_serial_tl_bits_out_bits_18_oe;
	wire iocell_serial_tl_bits_out_bits_19_pad;
	wire iocell_serial_tl_bits_out_bits_19_o;
	wire iocell_serial_tl_bits_out_bits_19_oe;
	wire iocell_serial_tl_bits_out_bits_20_pad;
	wire iocell_serial_tl_bits_out_bits_20_o;
	wire iocell_serial_tl_bits_out_bits_20_oe;
	wire iocell_serial_tl_bits_out_bits_21_pad;
	wire iocell_serial_tl_bits_out_bits_21_o;
	wire iocell_serial_tl_bits_out_bits_21_oe;
	wire iocell_serial_tl_bits_out_bits_22_pad;
	wire iocell_serial_tl_bits_out_bits_22_o;
	wire iocell_serial_tl_bits_out_bits_22_oe;
	wire iocell_serial_tl_bits_out_bits_23_pad;
	wire iocell_serial_tl_bits_out_bits_23_o;
	wire iocell_serial_tl_bits_out_bits_23_oe;
	wire iocell_serial_tl_bits_out_bits_24_pad;
	wire iocell_serial_tl_bits_out_bits_24_o;
	wire iocell_serial_tl_bits_out_bits_24_oe;
	wire iocell_serial_tl_bits_out_bits_25_pad;
	wire iocell_serial_tl_bits_out_bits_25_o;
	wire iocell_serial_tl_bits_out_bits_25_oe;
	wire iocell_serial_tl_bits_out_bits_26_pad;
	wire iocell_serial_tl_bits_out_bits_26_o;
	wire iocell_serial_tl_bits_out_bits_26_oe;
	wire iocell_serial_tl_bits_out_bits_27_pad;
	wire iocell_serial_tl_bits_out_bits_27_o;
	wire iocell_serial_tl_bits_out_bits_27_oe;
	wire iocell_serial_tl_bits_out_bits_28_pad;
	wire iocell_serial_tl_bits_out_bits_28_o;
	wire iocell_serial_tl_bits_out_bits_28_oe;
	wire iocell_serial_tl_bits_out_bits_29_pad;
	wire iocell_serial_tl_bits_out_bits_29_o;
	wire iocell_serial_tl_bits_out_bits_29_oe;
	wire iocell_serial_tl_bits_out_bits_30_pad;
	wire iocell_serial_tl_bits_out_bits_30_o;
	wire iocell_serial_tl_bits_out_bits_30_oe;
	wire iocell_serial_tl_bits_out_bits_31_pad;
	wire iocell_serial_tl_bits_out_bits_31_o;
	wire iocell_serial_tl_bits_out_bits_31_oe;
	wire iocell_serial_tl_bits_out_valid_pad;
	wire iocell_serial_tl_bits_out_valid_o;
	wire iocell_serial_tl_bits_out_valid_oe;
	wire iocell_serial_tl_bits_out_ready_pad;
	wire iocell_serial_tl_bits_out_ready_i;
	wire iocell_serial_tl_bits_out_ready_ie;
	wire iocell_serial_tl_bits_in_bits_pad;
	wire iocell_serial_tl_bits_in_bits_i;
	wire iocell_serial_tl_bits_in_bits_ie;
	wire iocell_serial_tl_bits_in_bits_1_pad;
	wire iocell_serial_tl_bits_in_bits_1_i;
	wire iocell_serial_tl_bits_in_bits_1_ie;
	wire iocell_serial_tl_bits_in_bits_2_pad;
	wire iocell_serial_tl_bits_in_bits_2_i;
	wire iocell_serial_tl_bits_in_bits_2_ie;
	wire iocell_serial_tl_bits_in_bits_3_pad;
	wire iocell_serial_tl_bits_in_bits_3_i;
	wire iocell_serial_tl_bits_in_bits_3_ie;
	wire iocell_serial_tl_bits_in_bits_4_pad;
	wire iocell_serial_tl_bits_in_bits_4_i;
	wire iocell_serial_tl_bits_in_bits_4_ie;
	wire iocell_serial_tl_bits_in_bits_5_pad;
	wire iocell_serial_tl_bits_in_bits_5_i;
	wire iocell_serial_tl_bits_in_bits_5_ie;
	wire iocell_serial_tl_bits_in_bits_6_pad;
	wire iocell_serial_tl_bits_in_bits_6_i;
	wire iocell_serial_tl_bits_in_bits_6_ie;
	wire iocell_serial_tl_bits_in_bits_7_pad;
	wire iocell_serial_tl_bits_in_bits_7_i;
	wire iocell_serial_tl_bits_in_bits_7_ie;
	wire iocell_serial_tl_bits_in_bits_8_pad;
	wire iocell_serial_tl_bits_in_bits_8_i;
	wire iocell_serial_tl_bits_in_bits_8_ie;
	wire iocell_serial_tl_bits_in_bits_9_pad;
	wire iocell_serial_tl_bits_in_bits_9_i;
	wire iocell_serial_tl_bits_in_bits_9_ie;
	wire iocell_serial_tl_bits_in_bits_10_pad;
	wire iocell_serial_tl_bits_in_bits_10_i;
	wire iocell_serial_tl_bits_in_bits_10_ie;
	wire iocell_serial_tl_bits_in_bits_11_pad;
	wire iocell_serial_tl_bits_in_bits_11_i;
	wire iocell_serial_tl_bits_in_bits_11_ie;
	wire iocell_serial_tl_bits_in_bits_12_pad;
	wire iocell_serial_tl_bits_in_bits_12_i;
	wire iocell_serial_tl_bits_in_bits_12_ie;
	wire iocell_serial_tl_bits_in_bits_13_pad;
	wire iocell_serial_tl_bits_in_bits_13_i;
	wire iocell_serial_tl_bits_in_bits_13_ie;
	wire iocell_serial_tl_bits_in_bits_14_pad;
	wire iocell_serial_tl_bits_in_bits_14_i;
	wire iocell_serial_tl_bits_in_bits_14_ie;
	wire iocell_serial_tl_bits_in_bits_15_pad;
	wire iocell_serial_tl_bits_in_bits_15_i;
	wire iocell_serial_tl_bits_in_bits_15_ie;
	wire iocell_serial_tl_bits_in_bits_16_pad;
	wire iocell_serial_tl_bits_in_bits_16_i;
	wire iocell_serial_tl_bits_in_bits_16_ie;
	wire iocell_serial_tl_bits_in_bits_17_pad;
	wire iocell_serial_tl_bits_in_bits_17_i;
	wire iocell_serial_tl_bits_in_bits_17_ie;
	wire iocell_serial_tl_bits_in_bits_18_pad;
	wire iocell_serial_tl_bits_in_bits_18_i;
	wire iocell_serial_tl_bits_in_bits_18_ie;
	wire iocell_serial_tl_bits_in_bits_19_pad;
	wire iocell_serial_tl_bits_in_bits_19_i;
	wire iocell_serial_tl_bits_in_bits_19_ie;
	wire iocell_serial_tl_bits_in_bits_20_pad;
	wire iocell_serial_tl_bits_in_bits_20_i;
	wire iocell_serial_tl_bits_in_bits_20_ie;
	wire iocell_serial_tl_bits_in_bits_21_pad;
	wire iocell_serial_tl_bits_in_bits_21_i;
	wire iocell_serial_tl_bits_in_bits_21_ie;
	wire iocell_serial_tl_bits_in_bits_22_pad;
	wire iocell_serial_tl_bits_in_bits_22_i;
	wire iocell_serial_tl_bits_in_bits_22_ie;
	wire iocell_serial_tl_bits_in_bits_23_pad;
	wire iocell_serial_tl_bits_in_bits_23_i;
	wire iocell_serial_tl_bits_in_bits_23_ie;
	wire iocell_serial_tl_bits_in_bits_24_pad;
	wire iocell_serial_tl_bits_in_bits_24_i;
	wire iocell_serial_tl_bits_in_bits_24_ie;
	wire iocell_serial_tl_bits_in_bits_25_pad;
	wire iocell_serial_tl_bits_in_bits_25_i;
	wire iocell_serial_tl_bits_in_bits_25_ie;
	wire iocell_serial_tl_bits_in_bits_26_pad;
	wire iocell_serial_tl_bits_in_bits_26_i;
	wire iocell_serial_tl_bits_in_bits_26_ie;
	wire iocell_serial_tl_bits_in_bits_27_pad;
	wire iocell_serial_tl_bits_in_bits_27_i;
	wire iocell_serial_tl_bits_in_bits_27_ie;
	wire iocell_serial_tl_bits_in_bits_28_pad;
	wire iocell_serial_tl_bits_in_bits_28_i;
	wire iocell_serial_tl_bits_in_bits_28_ie;
	wire iocell_serial_tl_bits_in_bits_29_pad;
	wire iocell_serial_tl_bits_in_bits_29_i;
	wire iocell_serial_tl_bits_in_bits_29_ie;
	wire iocell_serial_tl_bits_in_bits_30_pad;
	wire iocell_serial_tl_bits_in_bits_30_i;
	wire iocell_serial_tl_bits_in_bits_30_ie;
	wire iocell_serial_tl_bits_in_bits_31_pad;
	wire iocell_serial_tl_bits_in_bits_31_i;
	wire iocell_serial_tl_bits_in_bits_31_ie;
	wire iocell_serial_tl_bits_in_valid_pad;
	wire iocell_serial_tl_bits_in_valid_i;
	wire iocell_serial_tl_bits_in_valid_ie;
	wire iocell_serial_tl_bits_in_ready_pad;
	wire iocell_serial_tl_bits_in_ready_o;
	wire iocell_serial_tl_bits_in_ready_oe;
	wire iocell_serial_tl_clock_pad;
	wire iocell_serial_tl_clock_o;
	wire iocell_serial_tl_clock_oe;
	wire iocell_custom_boot_pad;
	wire iocell_custom_boot_i;
	wire iocell_custom_boot_ie;
	wire iocell_clock_clock_pad;
	wire iocell_clock_clock_i;
	wire iocell_clock_clock_ie;
	wire iocell_reset_pad;
	wire iocell_reset_i;
	wire iocell_reset_ie;
	wire iocell_uart_0_rxd_pad;
	wire iocell_uart_0_rxd_i;
	wire iocell_uart_0_rxd_ie;
	wire iocell_uart_0_txd_pad;
	wire iocell_uart_0_txd_o;
	wire iocell_uart_0_txd_oe;
	wire _debug_reset_syncd_WIRE = debug_reset_syncd_debug_reset_sync_io_q;
	wire _T = ~_debug_reset_syncd_WIRE;
	wire bundleIn_0_clock = system_auto_subsystem_cbus_fixedClockNode_out_clock;
	reg clock_en;
	wire [7:0] serial_tl_bits_out_bits_lo_lo = {iocell_serial_tl_bits_out_bits_7_pad, iocell_serial_tl_bits_out_bits_6_pad, iocell_serial_tl_bits_out_bits_5_pad, iocell_serial_tl_bits_out_bits_4_pad, iocell_serial_tl_bits_out_bits_3_pad, iocell_serial_tl_bits_out_bits_2_pad, iocell_serial_tl_bits_out_bits_1_pad, iocell_serial_tl_bits_out_bits_pad};
	wire [15:0] serial_tl_bits_out_bits_lo = {iocell_serial_tl_bits_out_bits_15_pad, iocell_serial_tl_bits_out_bits_14_pad, iocell_serial_tl_bits_out_bits_13_pad, iocell_serial_tl_bits_out_bits_12_pad, iocell_serial_tl_bits_out_bits_11_pad, iocell_serial_tl_bits_out_bits_10_pad, iocell_serial_tl_bits_out_bits_9_pad, iocell_serial_tl_bits_out_bits_8_pad, serial_tl_bits_out_bits_lo_lo};
	wire [7:0] serial_tl_bits_out_bits_hi_lo = {iocell_serial_tl_bits_out_bits_23_pad, iocell_serial_tl_bits_out_bits_22_pad, iocell_serial_tl_bits_out_bits_21_pad, iocell_serial_tl_bits_out_bits_20_pad, iocell_serial_tl_bits_out_bits_19_pad, iocell_serial_tl_bits_out_bits_18_pad, iocell_serial_tl_bits_out_bits_17_pad, iocell_serial_tl_bits_out_bits_16_pad};
	wire [15:0] serial_tl_bits_out_bits_hi = {iocell_serial_tl_bits_out_bits_31_pad, iocell_serial_tl_bits_out_bits_30_pad, iocell_serial_tl_bits_out_bits_29_pad, iocell_serial_tl_bits_out_bits_28_pad, iocell_serial_tl_bits_out_bits_27_pad, iocell_serial_tl_bits_out_bits_26_pad, iocell_serial_tl_bits_out_bits_25_pad, iocell_serial_tl_bits_out_bits_24_pad, serial_tl_bits_out_bits_hi_lo};
	wire [7:0] system_serial_tl_bits_in_bits_lo_lo = {iocell_serial_tl_bits_in_bits_7_i, iocell_serial_tl_bits_in_bits_6_i, iocell_serial_tl_bits_in_bits_5_i, iocell_serial_tl_bits_in_bits_4_i, iocell_serial_tl_bits_in_bits_3_i, iocell_serial_tl_bits_in_bits_2_i, iocell_serial_tl_bits_in_bits_1_i, iocell_serial_tl_bits_in_bits_i};
	wire [15:0] system_serial_tl_bits_in_bits_lo = {iocell_serial_tl_bits_in_bits_15_i, iocell_serial_tl_bits_in_bits_14_i, iocell_serial_tl_bits_in_bits_13_i, iocell_serial_tl_bits_in_bits_12_i, iocell_serial_tl_bits_in_bits_11_i, iocell_serial_tl_bits_in_bits_10_i, iocell_serial_tl_bits_in_bits_9_i, iocell_serial_tl_bits_in_bits_8_i, system_serial_tl_bits_in_bits_lo_lo};
	wire [7:0] system_serial_tl_bits_in_bits_hi_lo = {iocell_serial_tl_bits_in_bits_23_i, iocell_serial_tl_bits_in_bits_22_i, iocell_serial_tl_bits_in_bits_21_i, iocell_serial_tl_bits_in_bits_20_i, iocell_serial_tl_bits_in_bits_19_i, iocell_serial_tl_bits_in_bits_18_i, iocell_serial_tl_bits_in_bits_17_i, iocell_serial_tl_bits_in_bits_16_i};
	wire [15:0] system_serial_tl_bits_in_bits_hi = {iocell_serial_tl_bits_in_bits_31_i, iocell_serial_tl_bits_in_bits_30_i, iocell_serial_tl_bits_in_bits_29_i, iocell_serial_tl_bits_in_bits_28_i, iocell_serial_tl_bits_in_bits_27_i, iocell_serial_tl_bits_in_bits_26_i, iocell_serial_tl_bits_in_bits_25_i, iocell_serial_tl_bits_in_bits_24_i, system_serial_tl_bits_in_bits_hi_lo};
	DigitalTop system(
		.clock(system_clock),
		.reset(system_reset),
		.auto_implicitClockGrouper_out_clock(system_auto_implicitClockGrouper_out_clock),
		.auto_implicitClockGrouper_out_reset(system_auto_implicitClockGrouper_out_reset),
		.auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock(system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock),
		.auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset(system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset),
		.auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock(system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock),
		.auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset(system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset),
		.auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock(system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock),
		.auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset(system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset),
		.auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock(system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock),
		.auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset(system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset),
		.auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock(system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock),
		.auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset(system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset),
		.auto_subsystem_cbus_fixedClockNode_out_clock(system_auto_subsystem_cbus_fixedClockNode_out_clock),
		.auto_subsystem_cbus_fixedClockNode_out_reset(system_auto_subsystem_cbus_fixedClockNode_out_reset),
		.custom_boot(system_custom_boot),
		.serial_tl_clock(system_serial_tl_clock),
		.serial_tl_bits_in_ready(system_serial_tl_bits_in_ready),
		.serial_tl_bits_in_valid(system_serial_tl_bits_in_valid),
		.serial_tl_bits_in_bits(system_serial_tl_bits_in_bits),
		.serial_tl_bits_out_ready(system_serial_tl_bits_out_ready),
		.serial_tl_bits_out_valid(system_serial_tl_bits_out_valid),
		.serial_tl_bits_out_bits(system_serial_tl_bits_out_bits),
		.resetctrl_hartIsInReset_0(system_resetctrl_hartIsInReset_0),
		.debug_clock(system_debug_clock),
		.debug_reset(system_debug_reset),
		.debug_systemjtag_jtag_TCK(system_debug_systemjtag_jtag_TCK),
		.debug_systemjtag_jtag_TMS(system_debug_systemjtag_jtag_TMS),
		.debug_systemjtag_jtag_TDI(system_debug_systemjtag_jtag_TDI),
		.debug_systemjtag_jtag_TDO_data(system_debug_systemjtag_jtag_TDO_data),
		.debug_systemjtag_reset(system_debug_systemjtag_reset),
		.debug_dmactive(system_debug_dmactive),
		.debug_dmactiveAck(system_debug_dmactiveAck),
		.uart_0_txd(system_uart_0_txd),
		.uart_0_rxd(system_uart_0_rxd)
	);
	DividerOnlyClockGenerator dividerOnlyClockGen(
		.auto_divider_only_clock_gen_in_clock(dividerOnlyClockGen_auto_divider_only_clock_gen_in_clock),
		.auto_divider_only_clock_gen_in_reset(dividerOnlyClockGen_auto_divider_only_clock_gen_in_reset),
		.auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_clock(dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_clock),
		.auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_reset(dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_reset),
		.auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_clock(dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_clock),
		.auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_reset(dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_reset),
		.auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_clock(dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_clock),
		.auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_reset(dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_reset),
		.auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_clock(dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_clock),
		.auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_reset(dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_reset),
		.auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_clock(dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_clock),
		.auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_reset(dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_reset)
	);
	ResetCatchAndSync_d3 system_debug_systemjtag_reset_catcher(
		.clock(system_debug_systemjtag_reset_catcher_clock),
		.reset(system_debug_systemjtag_reset_catcher_reset),
		.io_sync_reset(system_debug_systemjtag_reset_catcher_io_sync_reset)
	);
	AsyncResetSynchronizerShiftReg_w1_d3_i0 debug_reset_syncd_debug_reset_sync(
		.clock(debug_reset_syncd_debug_reset_sync_clock),
		.reset(debug_reset_syncd_debug_reset_sync_reset),
		.io_d(debug_reset_syncd_debug_reset_sync_io_d),
		.io_q(debug_reset_syncd_debug_reset_sync_io_q)
	);
	ResetSynchronizerShiftReg_w1_d3_i0 dmactiveAck_dmactiveAck(
		.clock(dmactiveAck_dmactiveAck_clock),
		.reset(dmactiveAck_dmactiveAck_reset),
		.io_d(dmactiveAck_dmactiveAck_io_d),
		.io_q(dmactiveAck_dmactiveAck_io_q)
	);
	EICG_wrapper gated_clock_debug_clock_gate(
		.in(gated_clock_debug_clock_gate_in),
		.test_en(gated_clock_debug_clock_gate_test_en),
		.en(gated_clock_debug_clock_gate_en),
		.out(gated_clock_debug_clock_gate_out)
	);
	GenericDigitalOutIOCell iocell_jtag_TDO(
		.pad(iocell_jtag_TDO_pad),
		.o(iocell_jtag_TDO_o),
		.oe(iocell_jtag_TDO_oe)
	);
	GenericDigitalInIOCell iocell_jtag_TDI(
		.pad(iocell_jtag_TDI_pad),
		.i(iocell_jtag_TDI_i),
		.ie(iocell_jtag_TDI_ie)
	);
	GenericDigitalInIOCell iocell_jtag_TMS(
		.pad(iocell_jtag_TMS_pad),
		.i(iocell_jtag_TMS_i),
		.ie(iocell_jtag_TMS_ie)
	);
	GenericDigitalInIOCell iocell_jtag_TCK(
		.pad(iocell_jtag_TCK_pad),
		.i(iocell_jtag_TCK_i),
		.ie(iocell_jtag_TCK_ie)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits(
		.pad(iocell_serial_tl_bits_out_bits_pad),
		.o(iocell_serial_tl_bits_out_bits_o),
		.oe(iocell_serial_tl_bits_out_bits_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_1(
		.pad(iocell_serial_tl_bits_out_bits_1_pad),
		.o(iocell_serial_tl_bits_out_bits_1_o),
		.oe(iocell_serial_tl_bits_out_bits_1_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_2(
		.pad(iocell_serial_tl_bits_out_bits_2_pad),
		.o(iocell_serial_tl_bits_out_bits_2_o),
		.oe(iocell_serial_tl_bits_out_bits_2_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_3(
		.pad(iocell_serial_tl_bits_out_bits_3_pad),
		.o(iocell_serial_tl_bits_out_bits_3_o),
		.oe(iocell_serial_tl_bits_out_bits_3_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_4(
		.pad(iocell_serial_tl_bits_out_bits_4_pad),
		.o(iocell_serial_tl_bits_out_bits_4_o),
		.oe(iocell_serial_tl_bits_out_bits_4_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_5(
		.pad(iocell_serial_tl_bits_out_bits_5_pad),
		.o(iocell_serial_tl_bits_out_bits_5_o),
		.oe(iocell_serial_tl_bits_out_bits_5_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_6(
		.pad(iocell_serial_tl_bits_out_bits_6_pad),
		.o(iocell_serial_tl_bits_out_bits_6_o),
		.oe(iocell_serial_tl_bits_out_bits_6_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_7(
		.pad(iocell_serial_tl_bits_out_bits_7_pad),
		.o(iocell_serial_tl_bits_out_bits_7_o),
		.oe(iocell_serial_tl_bits_out_bits_7_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_8(
		.pad(iocell_serial_tl_bits_out_bits_8_pad),
		.o(iocell_serial_tl_bits_out_bits_8_o),
		.oe(iocell_serial_tl_bits_out_bits_8_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_9(
		.pad(iocell_serial_tl_bits_out_bits_9_pad),
		.o(iocell_serial_tl_bits_out_bits_9_o),
		.oe(iocell_serial_tl_bits_out_bits_9_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_10(
		.pad(iocell_serial_tl_bits_out_bits_10_pad),
		.o(iocell_serial_tl_bits_out_bits_10_o),
		.oe(iocell_serial_tl_bits_out_bits_10_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_11(
		.pad(iocell_serial_tl_bits_out_bits_11_pad),
		.o(iocell_serial_tl_bits_out_bits_11_o),
		.oe(iocell_serial_tl_bits_out_bits_11_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_12(
		.pad(iocell_serial_tl_bits_out_bits_12_pad),
		.o(iocell_serial_tl_bits_out_bits_12_o),
		.oe(iocell_serial_tl_bits_out_bits_12_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_13(
		.pad(iocell_serial_tl_bits_out_bits_13_pad),
		.o(iocell_serial_tl_bits_out_bits_13_o),
		.oe(iocell_serial_tl_bits_out_bits_13_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_14(
		.pad(iocell_serial_tl_bits_out_bits_14_pad),
		.o(iocell_serial_tl_bits_out_bits_14_o),
		.oe(iocell_serial_tl_bits_out_bits_14_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_15(
		.pad(iocell_serial_tl_bits_out_bits_15_pad),
		.o(iocell_serial_tl_bits_out_bits_15_o),
		.oe(iocell_serial_tl_bits_out_bits_15_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_16(
		.pad(iocell_serial_tl_bits_out_bits_16_pad),
		.o(iocell_serial_tl_bits_out_bits_16_o),
		.oe(iocell_serial_tl_bits_out_bits_16_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_17(
		.pad(iocell_serial_tl_bits_out_bits_17_pad),
		.o(iocell_serial_tl_bits_out_bits_17_o),
		.oe(iocell_serial_tl_bits_out_bits_17_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_18(
		.pad(iocell_serial_tl_bits_out_bits_18_pad),
		.o(iocell_serial_tl_bits_out_bits_18_o),
		.oe(iocell_serial_tl_bits_out_bits_18_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_19(
		.pad(iocell_serial_tl_bits_out_bits_19_pad),
		.o(iocell_serial_tl_bits_out_bits_19_o),
		.oe(iocell_serial_tl_bits_out_bits_19_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_20(
		.pad(iocell_serial_tl_bits_out_bits_20_pad),
		.o(iocell_serial_tl_bits_out_bits_20_o),
		.oe(iocell_serial_tl_bits_out_bits_20_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_21(
		.pad(iocell_serial_tl_bits_out_bits_21_pad),
		.o(iocell_serial_tl_bits_out_bits_21_o),
		.oe(iocell_serial_tl_bits_out_bits_21_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_22(
		.pad(iocell_serial_tl_bits_out_bits_22_pad),
		.o(iocell_serial_tl_bits_out_bits_22_o),
		.oe(iocell_serial_tl_bits_out_bits_22_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_23(
		.pad(iocell_serial_tl_bits_out_bits_23_pad),
		.o(iocell_serial_tl_bits_out_bits_23_o),
		.oe(iocell_serial_tl_bits_out_bits_23_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_24(
		.pad(iocell_serial_tl_bits_out_bits_24_pad),
		.o(iocell_serial_tl_bits_out_bits_24_o),
		.oe(iocell_serial_tl_bits_out_bits_24_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_25(
		.pad(iocell_serial_tl_bits_out_bits_25_pad),
		.o(iocell_serial_tl_bits_out_bits_25_o),
		.oe(iocell_serial_tl_bits_out_bits_25_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_26(
		.pad(iocell_serial_tl_bits_out_bits_26_pad),
		.o(iocell_serial_tl_bits_out_bits_26_o),
		.oe(iocell_serial_tl_bits_out_bits_26_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_27(
		.pad(iocell_serial_tl_bits_out_bits_27_pad),
		.o(iocell_serial_tl_bits_out_bits_27_o),
		.oe(iocell_serial_tl_bits_out_bits_27_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_28(
		.pad(iocell_serial_tl_bits_out_bits_28_pad),
		.o(iocell_serial_tl_bits_out_bits_28_o),
		.oe(iocell_serial_tl_bits_out_bits_28_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_29(
		.pad(iocell_serial_tl_bits_out_bits_29_pad),
		.o(iocell_serial_tl_bits_out_bits_29_o),
		.oe(iocell_serial_tl_bits_out_bits_29_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_30(
		.pad(iocell_serial_tl_bits_out_bits_30_pad),
		.o(iocell_serial_tl_bits_out_bits_30_o),
		.oe(iocell_serial_tl_bits_out_bits_30_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_bits_31(
		.pad(iocell_serial_tl_bits_out_bits_31_pad),
		.o(iocell_serial_tl_bits_out_bits_31_o),
		.oe(iocell_serial_tl_bits_out_bits_31_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_out_valid(
		.pad(iocell_serial_tl_bits_out_valid_pad),
		.o(iocell_serial_tl_bits_out_valid_o),
		.oe(iocell_serial_tl_bits_out_valid_oe)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_out_ready(
		.pad(iocell_serial_tl_bits_out_ready_pad),
		.i(iocell_serial_tl_bits_out_ready_i),
		.ie(iocell_serial_tl_bits_out_ready_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits(
		.pad(iocell_serial_tl_bits_in_bits_pad),
		.i(iocell_serial_tl_bits_in_bits_i),
		.ie(iocell_serial_tl_bits_in_bits_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_1(
		.pad(iocell_serial_tl_bits_in_bits_1_pad),
		.i(iocell_serial_tl_bits_in_bits_1_i),
		.ie(iocell_serial_tl_bits_in_bits_1_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_2(
		.pad(iocell_serial_tl_bits_in_bits_2_pad),
		.i(iocell_serial_tl_bits_in_bits_2_i),
		.ie(iocell_serial_tl_bits_in_bits_2_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_3(
		.pad(iocell_serial_tl_bits_in_bits_3_pad),
		.i(iocell_serial_tl_bits_in_bits_3_i),
		.ie(iocell_serial_tl_bits_in_bits_3_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_4(
		.pad(iocell_serial_tl_bits_in_bits_4_pad),
		.i(iocell_serial_tl_bits_in_bits_4_i),
		.ie(iocell_serial_tl_bits_in_bits_4_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_5(
		.pad(iocell_serial_tl_bits_in_bits_5_pad),
		.i(iocell_serial_tl_bits_in_bits_5_i),
		.ie(iocell_serial_tl_bits_in_bits_5_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_6(
		.pad(iocell_serial_tl_bits_in_bits_6_pad),
		.i(iocell_serial_tl_bits_in_bits_6_i),
		.ie(iocell_serial_tl_bits_in_bits_6_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_7(
		.pad(iocell_serial_tl_bits_in_bits_7_pad),
		.i(iocell_serial_tl_bits_in_bits_7_i),
		.ie(iocell_serial_tl_bits_in_bits_7_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_8(
		.pad(iocell_serial_tl_bits_in_bits_8_pad),
		.i(iocell_serial_tl_bits_in_bits_8_i),
		.ie(iocell_serial_tl_bits_in_bits_8_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_9(
		.pad(iocell_serial_tl_bits_in_bits_9_pad),
		.i(iocell_serial_tl_bits_in_bits_9_i),
		.ie(iocell_serial_tl_bits_in_bits_9_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_10(
		.pad(iocell_serial_tl_bits_in_bits_10_pad),
		.i(iocell_serial_tl_bits_in_bits_10_i),
		.ie(iocell_serial_tl_bits_in_bits_10_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_11(
		.pad(iocell_serial_tl_bits_in_bits_11_pad),
		.i(iocell_serial_tl_bits_in_bits_11_i),
		.ie(iocell_serial_tl_bits_in_bits_11_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_12(
		.pad(iocell_serial_tl_bits_in_bits_12_pad),
		.i(iocell_serial_tl_bits_in_bits_12_i),
		.ie(iocell_serial_tl_bits_in_bits_12_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_13(
		.pad(iocell_serial_tl_bits_in_bits_13_pad),
		.i(iocell_serial_tl_bits_in_bits_13_i),
		.ie(iocell_serial_tl_bits_in_bits_13_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_14(
		.pad(iocell_serial_tl_bits_in_bits_14_pad),
		.i(iocell_serial_tl_bits_in_bits_14_i),
		.ie(iocell_serial_tl_bits_in_bits_14_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_15(
		.pad(iocell_serial_tl_bits_in_bits_15_pad),
		.i(iocell_serial_tl_bits_in_bits_15_i),
		.ie(iocell_serial_tl_bits_in_bits_15_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_16(
		.pad(iocell_serial_tl_bits_in_bits_16_pad),
		.i(iocell_serial_tl_bits_in_bits_16_i),
		.ie(iocell_serial_tl_bits_in_bits_16_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_17(
		.pad(iocell_serial_tl_bits_in_bits_17_pad),
		.i(iocell_serial_tl_bits_in_bits_17_i),
		.ie(iocell_serial_tl_bits_in_bits_17_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_18(
		.pad(iocell_serial_tl_bits_in_bits_18_pad),
		.i(iocell_serial_tl_bits_in_bits_18_i),
		.ie(iocell_serial_tl_bits_in_bits_18_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_19(
		.pad(iocell_serial_tl_bits_in_bits_19_pad),
		.i(iocell_serial_tl_bits_in_bits_19_i),
		.ie(iocell_serial_tl_bits_in_bits_19_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_20(
		.pad(iocell_serial_tl_bits_in_bits_20_pad),
		.i(iocell_serial_tl_bits_in_bits_20_i),
		.ie(iocell_serial_tl_bits_in_bits_20_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_21(
		.pad(iocell_serial_tl_bits_in_bits_21_pad),
		.i(iocell_serial_tl_bits_in_bits_21_i),
		.ie(iocell_serial_tl_bits_in_bits_21_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_22(
		.pad(iocell_serial_tl_bits_in_bits_22_pad),
		.i(iocell_serial_tl_bits_in_bits_22_i),
		.ie(iocell_serial_tl_bits_in_bits_22_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_23(
		.pad(iocell_serial_tl_bits_in_bits_23_pad),
		.i(iocell_serial_tl_bits_in_bits_23_i),
		.ie(iocell_serial_tl_bits_in_bits_23_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_24(
		.pad(iocell_serial_tl_bits_in_bits_24_pad),
		.i(iocell_serial_tl_bits_in_bits_24_i),
		.ie(iocell_serial_tl_bits_in_bits_24_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_25(
		.pad(iocell_serial_tl_bits_in_bits_25_pad),
		.i(iocell_serial_tl_bits_in_bits_25_i),
		.ie(iocell_serial_tl_bits_in_bits_25_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_26(
		.pad(iocell_serial_tl_bits_in_bits_26_pad),
		.i(iocell_serial_tl_bits_in_bits_26_i),
		.ie(iocell_serial_tl_bits_in_bits_26_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_27(
		.pad(iocell_serial_tl_bits_in_bits_27_pad),
		.i(iocell_serial_tl_bits_in_bits_27_i),
		.ie(iocell_serial_tl_bits_in_bits_27_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_28(
		.pad(iocell_serial_tl_bits_in_bits_28_pad),
		.i(iocell_serial_tl_bits_in_bits_28_i),
		.ie(iocell_serial_tl_bits_in_bits_28_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_29(
		.pad(iocell_serial_tl_bits_in_bits_29_pad),
		.i(iocell_serial_tl_bits_in_bits_29_i),
		.ie(iocell_serial_tl_bits_in_bits_29_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_30(
		.pad(iocell_serial_tl_bits_in_bits_30_pad),
		.i(iocell_serial_tl_bits_in_bits_30_i),
		.ie(iocell_serial_tl_bits_in_bits_30_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_bits_31(
		.pad(iocell_serial_tl_bits_in_bits_31_pad),
		.i(iocell_serial_tl_bits_in_bits_31_i),
		.ie(iocell_serial_tl_bits_in_bits_31_ie)
	);
	GenericDigitalInIOCell iocell_serial_tl_bits_in_valid(
		.pad(iocell_serial_tl_bits_in_valid_pad),
		.i(iocell_serial_tl_bits_in_valid_i),
		.ie(iocell_serial_tl_bits_in_valid_ie)
	);
	GenericDigitalOutIOCell iocell_serial_tl_bits_in_ready(
		.pad(iocell_serial_tl_bits_in_ready_pad),
		.o(iocell_serial_tl_bits_in_ready_o),
		.oe(iocell_serial_tl_bits_in_ready_oe)
	);
	GenericDigitalOutIOCell iocell_serial_tl_clock(
		.pad(iocell_serial_tl_clock_pad),
		.o(iocell_serial_tl_clock_o),
		.oe(iocell_serial_tl_clock_oe)
	);
	GenericDigitalInIOCell iocell_custom_boot(
		.pad(iocell_custom_boot_pad),
		.i(iocell_custom_boot_i),
		.ie(iocell_custom_boot_ie)
	);
	GenericDigitalInIOCell iocell_clock_clock(
		.pad(iocell_clock_clock_pad),
		.i(iocell_clock_clock_i),
		.ie(iocell_clock_clock_ie)
	);
	GenericDigitalInIOCell iocell_reset(
		.pad(iocell_reset_pad),
		.i(iocell_reset_i),
		.ie(iocell_reset_ie)
	);
	GenericDigitalInIOCell iocell_uart_0_rxd(
		.pad(iocell_uart_0_rxd_pad),
		.i(iocell_uart_0_rxd_i),
		.ie(iocell_uart_0_rxd_ie)
	);
	GenericDigitalOutIOCell iocell_uart_0_txd(
		.pad(iocell_uart_0_txd_pad),
		.o(iocell_uart_0_txd_o),
		.oe(iocell_uart_0_txd_oe)
	);
	assign jtag_TDO = iocell_jtag_TDO_pad;
	assign serial_tl_clock = iocell_serial_tl_clock_pad;
	assign serial_tl_bits_in_ready = iocell_serial_tl_bits_in_ready_pad;
	assign serial_tl_bits_out_valid = iocell_serial_tl_bits_out_valid_pad;
	assign serial_tl_bits_out_bits = {serial_tl_bits_out_bits_hi, serial_tl_bits_out_bits_lo};
	assign uart_0_txd = iocell_uart_0_txd_pad;
	assign system_clock = system_auto_implicitClockGrouper_out_clock;
	assign system_reset = system_auto_implicitClockGrouper_out_reset;
	assign system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_clock = dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_clock;
	assign system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_implicit_clock_reset = dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_implicit_clock_reset;
	assign system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_clock = dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_clock;
	assign system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_cbus_0_reset = dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_cbus_0_reset;
	assign system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_clock = dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_clock;
	assign system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_fbus_0_reset = dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_fbus_0_reset;
	assign system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_clock = dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_clock;
	assign system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_pbus_0_reset = dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_pbus_0_reset;
	assign system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_clock = dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_clock;
	assign system_auto_prci_ctrl_domain_tileResetSetter_clock_in_member_allClocks_subsystem_sbus_0_reset = dividerOnlyClockGen_auto_divider_only_clock_gen_out_member_allClocks_subsystem_sbus_0_reset;
	assign system_custom_boot = iocell_custom_boot_i;
	assign system_serial_tl_bits_in_valid = iocell_serial_tl_bits_in_valid_i;
	assign system_serial_tl_bits_in_bits = {system_serial_tl_bits_in_bits_hi, system_serial_tl_bits_in_bits_lo};
	assign system_serial_tl_bits_out_ready = iocell_serial_tl_bits_out_ready_i;
	assign system_resetctrl_hartIsInReset_0 = system_auto_subsystem_cbus_fixedClockNode_out_reset;
	assign system_debug_clock = gated_clock_debug_clock_gate_out;
	assign system_debug_reset = ~_debug_reset_syncd_WIRE;
	assign system_debug_systemjtag_jtag_TCK = iocell_jtag_TCK_i;
	assign system_debug_systemjtag_jtag_TMS = iocell_jtag_TMS_i;
	assign system_debug_systemjtag_jtag_TDI = iocell_jtag_TDI_i;
	assign system_debug_systemjtag_reset = system_debug_systemjtag_reset_catcher_io_sync_reset;
	assign system_debug_dmactiveAck = dmactiveAck_dmactiveAck_io_q;
	assign system_uart_0_rxd = iocell_uart_0_rxd_i;
	assign dividerOnlyClockGen_auto_divider_only_clock_gen_in_clock = iocell_clock_clock_i;
	assign dividerOnlyClockGen_auto_divider_only_clock_gen_in_reset = iocell_reset_i;
	assign system_debug_systemjtag_reset_catcher_clock = system_debug_systemjtag_jtag_TCK;
	assign system_debug_systemjtag_reset_catcher_reset = system_auto_subsystem_cbus_fixedClockNode_out_reset;
	assign debug_reset_syncd_debug_reset_sync_clock = system_auto_subsystem_cbus_fixedClockNode_out_clock;
	assign debug_reset_syncd_debug_reset_sync_reset = system_debug_systemjtag_reset;
	assign debug_reset_syncd_debug_reset_sync_io_d = 1'h1;
	assign dmactiveAck_dmactiveAck_clock = system_auto_subsystem_cbus_fixedClockNode_out_clock;
	assign dmactiveAck_dmactiveAck_reset = ~_debug_reset_syncd_WIRE;
	assign dmactiveAck_dmactiveAck_io_d = system_debug_dmactive;
	assign gated_clock_debug_clock_gate_in = system_auto_subsystem_cbus_fixedClockNode_out_clock;
	assign gated_clock_debug_clock_gate_test_en = 1'h0;
	assign gated_clock_debug_clock_gate_en = clock_en;
	assign iocell_jtag_TDO_o = system_debug_systemjtag_jtag_TDO_data;
	assign iocell_jtag_TDO_oe = 1'h1;
	assign iocell_jtag_TDI_pad = jtag_TDI;
	assign iocell_jtag_TDI_ie = 1'h1;
	assign iocell_jtag_TMS_pad = jtag_TMS;
	assign iocell_jtag_TMS_ie = 1'h1;
	assign iocell_jtag_TCK_pad = jtag_TCK;
	assign iocell_jtag_TCK_ie = 1'h1;
	assign iocell_serial_tl_bits_out_bits_o = system_serial_tl_bits_out_bits[0];
	assign iocell_serial_tl_bits_out_bits_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_1_o = system_serial_tl_bits_out_bits[1];
	assign iocell_serial_tl_bits_out_bits_1_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_2_o = system_serial_tl_bits_out_bits[2];
	assign iocell_serial_tl_bits_out_bits_2_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_3_o = system_serial_tl_bits_out_bits[3];
	assign iocell_serial_tl_bits_out_bits_3_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_4_o = system_serial_tl_bits_out_bits[4];
	assign iocell_serial_tl_bits_out_bits_4_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_5_o = system_serial_tl_bits_out_bits[5];
	assign iocell_serial_tl_bits_out_bits_5_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_6_o = system_serial_tl_bits_out_bits[6];
	assign iocell_serial_tl_bits_out_bits_6_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_7_o = system_serial_tl_bits_out_bits[7];
	assign iocell_serial_tl_bits_out_bits_7_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_8_o = system_serial_tl_bits_out_bits[8];
	assign iocell_serial_tl_bits_out_bits_8_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_9_o = system_serial_tl_bits_out_bits[9];
	assign iocell_serial_tl_bits_out_bits_9_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_10_o = system_serial_tl_bits_out_bits[10];
	assign iocell_serial_tl_bits_out_bits_10_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_11_o = system_serial_tl_bits_out_bits[11];
	assign iocell_serial_tl_bits_out_bits_11_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_12_o = system_serial_tl_bits_out_bits[12];
	assign iocell_serial_tl_bits_out_bits_12_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_13_o = system_serial_tl_bits_out_bits[13];
	assign iocell_serial_tl_bits_out_bits_13_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_14_o = system_serial_tl_bits_out_bits[14];
	assign iocell_serial_tl_bits_out_bits_14_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_15_o = system_serial_tl_bits_out_bits[15];
	assign iocell_serial_tl_bits_out_bits_15_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_16_o = system_serial_tl_bits_out_bits[16];
	assign iocell_serial_tl_bits_out_bits_16_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_17_o = system_serial_tl_bits_out_bits[17];
	assign iocell_serial_tl_bits_out_bits_17_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_18_o = system_serial_tl_bits_out_bits[18];
	assign iocell_serial_tl_bits_out_bits_18_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_19_o = system_serial_tl_bits_out_bits[19];
	assign iocell_serial_tl_bits_out_bits_19_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_20_o = system_serial_tl_bits_out_bits[20];
	assign iocell_serial_tl_bits_out_bits_20_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_21_o = system_serial_tl_bits_out_bits[21];
	assign iocell_serial_tl_bits_out_bits_21_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_22_o = system_serial_tl_bits_out_bits[22];
	assign iocell_serial_tl_bits_out_bits_22_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_23_o = system_serial_tl_bits_out_bits[23];
	assign iocell_serial_tl_bits_out_bits_23_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_24_o = system_serial_tl_bits_out_bits[24];
	assign iocell_serial_tl_bits_out_bits_24_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_25_o = system_serial_tl_bits_out_bits[25];
	assign iocell_serial_tl_bits_out_bits_25_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_26_o = system_serial_tl_bits_out_bits[26];
	assign iocell_serial_tl_bits_out_bits_26_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_27_o = system_serial_tl_bits_out_bits[27];
	assign iocell_serial_tl_bits_out_bits_27_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_28_o = system_serial_tl_bits_out_bits[28];
	assign iocell_serial_tl_bits_out_bits_28_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_29_o = system_serial_tl_bits_out_bits[29];
	assign iocell_serial_tl_bits_out_bits_29_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_30_o = system_serial_tl_bits_out_bits[30];
	assign iocell_serial_tl_bits_out_bits_30_oe = 1'h1;
	assign iocell_serial_tl_bits_out_bits_31_o = system_serial_tl_bits_out_bits[31];
	assign iocell_serial_tl_bits_out_bits_31_oe = 1'h1;
	assign iocell_serial_tl_bits_out_valid_o = system_serial_tl_bits_out_valid;
	assign iocell_serial_tl_bits_out_valid_oe = 1'h1;
	assign iocell_serial_tl_bits_out_ready_pad = serial_tl_bits_out_ready;
	assign iocell_serial_tl_bits_out_ready_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_pad = serial_tl_bits_in_bits[0];
	assign iocell_serial_tl_bits_in_bits_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_1_pad = serial_tl_bits_in_bits[1];
	assign iocell_serial_tl_bits_in_bits_1_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_2_pad = serial_tl_bits_in_bits[2];
	assign iocell_serial_tl_bits_in_bits_2_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_3_pad = serial_tl_bits_in_bits[3];
	assign iocell_serial_tl_bits_in_bits_3_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_4_pad = serial_tl_bits_in_bits[4];
	assign iocell_serial_tl_bits_in_bits_4_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_5_pad = serial_tl_bits_in_bits[5];
	assign iocell_serial_tl_bits_in_bits_5_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_6_pad = serial_tl_bits_in_bits[6];
	assign iocell_serial_tl_bits_in_bits_6_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_7_pad = serial_tl_bits_in_bits[7];
	assign iocell_serial_tl_bits_in_bits_7_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_8_pad = serial_tl_bits_in_bits[8];
	assign iocell_serial_tl_bits_in_bits_8_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_9_pad = serial_tl_bits_in_bits[9];
	assign iocell_serial_tl_bits_in_bits_9_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_10_pad = serial_tl_bits_in_bits[10];
	assign iocell_serial_tl_bits_in_bits_10_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_11_pad = serial_tl_bits_in_bits[11];
	assign iocell_serial_tl_bits_in_bits_11_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_12_pad = serial_tl_bits_in_bits[12];
	assign iocell_serial_tl_bits_in_bits_12_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_13_pad = serial_tl_bits_in_bits[13];
	assign iocell_serial_tl_bits_in_bits_13_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_14_pad = serial_tl_bits_in_bits[14];
	assign iocell_serial_tl_bits_in_bits_14_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_15_pad = serial_tl_bits_in_bits[15];
	assign iocell_serial_tl_bits_in_bits_15_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_16_pad = serial_tl_bits_in_bits[16];
	assign iocell_serial_tl_bits_in_bits_16_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_17_pad = serial_tl_bits_in_bits[17];
	assign iocell_serial_tl_bits_in_bits_17_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_18_pad = serial_tl_bits_in_bits[18];
	assign iocell_serial_tl_bits_in_bits_18_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_19_pad = serial_tl_bits_in_bits[19];
	assign iocell_serial_tl_bits_in_bits_19_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_20_pad = serial_tl_bits_in_bits[20];
	assign iocell_serial_tl_bits_in_bits_20_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_21_pad = serial_tl_bits_in_bits[21];
	assign iocell_serial_tl_bits_in_bits_21_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_22_pad = serial_tl_bits_in_bits[22];
	assign iocell_serial_tl_bits_in_bits_22_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_23_pad = serial_tl_bits_in_bits[23];
	assign iocell_serial_tl_bits_in_bits_23_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_24_pad = serial_tl_bits_in_bits[24];
	assign iocell_serial_tl_bits_in_bits_24_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_25_pad = serial_tl_bits_in_bits[25];
	assign iocell_serial_tl_bits_in_bits_25_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_26_pad = serial_tl_bits_in_bits[26];
	assign iocell_serial_tl_bits_in_bits_26_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_27_pad = serial_tl_bits_in_bits[27];
	assign iocell_serial_tl_bits_in_bits_27_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_28_pad = serial_tl_bits_in_bits[28];
	assign iocell_serial_tl_bits_in_bits_28_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_29_pad = serial_tl_bits_in_bits[29];
	assign iocell_serial_tl_bits_in_bits_29_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_30_pad = serial_tl_bits_in_bits[30];
	assign iocell_serial_tl_bits_in_bits_30_ie = 1'h1;
	assign iocell_serial_tl_bits_in_bits_31_pad = serial_tl_bits_in_bits[31];
	assign iocell_serial_tl_bits_in_bits_31_ie = 1'h1;
	assign iocell_serial_tl_bits_in_valid_pad = serial_tl_bits_in_valid;
	assign iocell_serial_tl_bits_in_valid_ie = 1'h1;
	assign iocell_serial_tl_bits_in_ready_o = system_serial_tl_bits_in_ready;
	assign iocell_serial_tl_bits_in_ready_oe = 1'h1;
	assign iocell_serial_tl_clock_o = system_serial_tl_clock;
	assign iocell_serial_tl_clock_oe = 1'h1;
	assign iocell_custom_boot_pad = custom_boot;
	assign iocell_custom_boot_ie = 1'h1;
	assign iocell_clock_clock_pad = clock_clock;
	assign iocell_clock_clock_ie = 1'h1;
	assign iocell_reset_pad = reset;
	assign iocell_reset_ie = 1'h1;
	assign iocell_uart_0_rxd_pad = uart_0_rxd;
	assign iocell_uart_0_rxd_ie = 1'h1;
	assign iocell_uart_0_txd_o = system_uart_0_txd;
	assign iocell_uart_0_txd_oe = 1'h1;
	always @(posedge bundleIn_0_clock or posedge _T)
		if (_T)
			clock_en <= 1'h1;
		else
			clock_en <= dmactiveAck_dmactiveAck_io_q;
endmodule
module data_arrays_0 (
	RW0_addr,
	RW0_en,
	RW0_clk,
	RW0_wmode,
	RW0_wdata_0,
	RW0_wdata_1,
	RW0_wdata_2,
	RW0_wdata_3,
	RW0_rdata_0,
	RW0_rdata_1,
	RW0_rdata_2,
	RW0_rdata_3,
	RW0_wmask_0,
	RW0_wmask_1,
	RW0_wmask_2,
	RW0_wmask_3
);
	input [11:0] RW0_addr;
	input RW0_en;
	input RW0_clk;
	input RW0_wmode;
	input [7:0] RW0_wdata_0;
	input [7:0] RW0_wdata_1;
	input [7:0] RW0_wdata_2;
	input [7:0] RW0_wdata_3;
	output wire [7:0] RW0_rdata_0;
	output wire [7:0] RW0_rdata_1;
	output wire [7:0] RW0_rdata_2;
	output wire [7:0] RW0_rdata_3;
	input RW0_wmask_0;
	input RW0_wmask_1;
	input RW0_wmask_2;
	input RW0_wmask_3;
	wire [11:0] data_arrays_0_ext_RW0_addr;
	wire data_arrays_0_ext_RW0_en;
	wire data_arrays_0_ext_RW0_clk;
	wire data_arrays_0_ext_RW0_wmode;
	wire [31:0] data_arrays_0_ext_RW0_wdata;
	wire [31:0] data_arrays_0_ext_RW0_rdata;
	wire [3:0] data_arrays_0_ext_RW0_wmask;
	wire [15:0] _GEN_0 = {RW0_wdata_3, RW0_wdata_2};
	wire [15:0] _GEN_1 = {RW0_wdata_1, RW0_wdata_0};
	wire [1:0] _GEN_2 = {RW0_wmask_3, RW0_wmask_2};
	wire [1:0] _GEN_3 = {RW0_wmask_1, RW0_wmask_0};
	data_arrays_0_ext data_arrays_0_ext(
		.RW0_addr(data_arrays_0_ext_RW0_addr),
		.RW0_en(data_arrays_0_ext_RW0_en),
		.RW0_clk(data_arrays_0_ext_RW0_clk),
		.RW0_wmode(data_arrays_0_ext_RW0_wmode),
		.RW0_wdata(data_arrays_0_ext_RW0_wdata),
		.RW0_rdata(data_arrays_0_ext_RW0_rdata),
		.RW0_wmask(data_arrays_0_ext_RW0_wmask)
	);
	assign data_arrays_0_ext_RW0_clk = RW0_clk;
	assign data_arrays_0_ext_RW0_en = RW0_en;
	assign data_arrays_0_ext_RW0_addr = RW0_addr;
	assign RW0_rdata_0 = data_arrays_0_ext_RW0_rdata[7:0];
	assign RW0_rdata_1 = data_arrays_0_ext_RW0_rdata[15:8];
	assign RW0_rdata_2 = data_arrays_0_ext_RW0_rdata[23:16];
	assign RW0_rdata_3 = data_arrays_0_ext_RW0_rdata[31:24];
	assign data_arrays_0_ext_RW0_wmode = RW0_wmode;
	assign data_arrays_0_ext_RW0_wdata = {_GEN_0, _GEN_1};
	assign data_arrays_0_ext_RW0_wmask = {_GEN_2, _GEN_3};
endmodule
module tag_array (
	RW0_addr,
	RW0_en,
	RW0_clk,
	RW0_wmode,
	RW0_wdata_0,
	RW0_rdata_0
);
	input [5:0] RW0_addr;
	input RW0_en;
	input RW0_clk;
	input RW0_wmode;
	input [20:0] RW0_wdata_0;
	output wire [20:0] RW0_rdata_0;
	wire [5:0] tag_array_ext_RW0_addr;
	wire tag_array_ext_RW0_en;
	wire tag_array_ext_RW0_clk;
	wire tag_array_ext_RW0_wmode;
	wire [20:0] tag_array_ext_RW0_wdata;
	wire [20:0] tag_array_ext_RW0_rdata;
	wire tag_array_ext_RW0_wmask;
	tag_array_ext tag_array_ext(
		.RW0_addr(tag_array_ext_RW0_addr),
		.RW0_en(tag_array_ext_RW0_en),
		.RW0_clk(tag_array_ext_RW0_clk),
		.RW0_wmode(tag_array_ext_RW0_wmode),
		.RW0_wdata(tag_array_ext_RW0_wdata),
		.RW0_rdata(tag_array_ext_RW0_rdata),
		.RW0_wmask(tag_array_ext_RW0_wmask)
	);
	assign tag_array_ext_RW0_clk = RW0_clk;
	assign tag_array_ext_RW0_en = RW0_en;
	assign tag_array_ext_RW0_addr = RW0_addr;
	assign RW0_rdata_0 = tag_array_ext_RW0_rdata;
	assign tag_array_ext_RW0_wmode = RW0_wmode;
	assign tag_array_ext_RW0_wdata = RW0_wdata_0;
	assign tag_array_ext_RW0_wmask = 1'h1;
endmodule
module data_arrays_0_0 (
	RW0_addr,
	RW0_en,
	RW0_clk,
	RW0_wmode,
	RW0_wdata_0,
	RW0_rdata_0
);
	input [9:0] RW0_addr;
	input RW0_en;
	input RW0_clk;
	input RW0_wmode;
	input [31:0] RW0_wdata_0;
	output wire [31:0] RW0_rdata_0;
	wire [9:0] data_arrays_0_0_ext_RW0_addr;
	wire data_arrays_0_0_ext_RW0_en;
	wire data_arrays_0_0_ext_RW0_clk;
	wire data_arrays_0_0_ext_RW0_wmode;
	wire [31:0] data_arrays_0_0_ext_RW0_wdata;
	wire [31:0] data_arrays_0_0_ext_RW0_rdata;
	wire data_arrays_0_0_ext_RW0_wmask;
	data_arrays_0_0_ext data_arrays_0_0_ext(
		.RW0_addr(data_arrays_0_0_ext_RW0_addr),
		.RW0_en(data_arrays_0_0_ext_RW0_en),
		.RW0_clk(data_arrays_0_0_ext_RW0_clk),
		.RW0_wmode(data_arrays_0_0_ext_RW0_wmode),
		.RW0_wdata(data_arrays_0_0_ext_RW0_wdata),
		.RW0_rdata(data_arrays_0_0_ext_RW0_rdata),
		.RW0_wmask(data_arrays_0_0_ext_RW0_wmask)
	);
	assign data_arrays_0_0_ext_RW0_clk = RW0_clk;
	assign data_arrays_0_0_ext_RW0_en = RW0_en;
	assign data_arrays_0_0_ext_RW0_addr = RW0_addr;
	assign RW0_rdata_0 = data_arrays_0_0_ext_RW0_rdata;
	assign data_arrays_0_0_ext_RW0_wmode = RW0_wmode;
	assign data_arrays_0_0_ext_RW0_wdata = RW0_wdata_0;
	assign data_arrays_0_0_ext_RW0_wmask = 1'h1;
endmodule
module l2_tlb_ram (
	RW0_clk,
	RW0_wdata_0
);
	input RW0_clk;
	input [36:0] RW0_wdata_0;
	wire [9:0] l2_tlb_ram_ext_RW0_addr;
	wire l2_tlb_ram_ext_RW0_en;
	wire l2_tlb_ram_ext_RW0_clk;
	wire l2_tlb_ram_ext_RW0_wmode;
	wire [36:0] l2_tlb_ram_ext_RW0_wdata;
	wire [36:0] l2_tlb_ram_ext_RW0_rdata;
	l2_tlb_ram_ext l2_tlb_ram_ext(
		.RW0_addr(l2_tlb_ram_ext_RW0_addr),
		.RW0_en(l2_tlb_ram_ext_RW0_en),
		.RW0_clk(l2_tlb_ram_ext_RW0_clk),
		.RW0_wmode(l2_tlb_ram_ext_RW0_wmode),
		.RW0_wdata(l2_tlb_ram_ext_RW0_wdata),
		.RW0_rdata(l2_tlb_ram_ext_RW0_rdata)
	);
	assign l2_tlb_ram_ext_RW0_clk = RW0_clk;
	assign l2_tlb_ram_ext_RW0_en = 1'h0;
	assign l2_tlb_ram_ext_RW0_addr = 10'h000;
	assign l2_tlb_ram_ext_RW0_wmode = 1'h0;
	assign l2_tlb_ram_ext_RW0_wdata = RW0_wdata_0;
endmodule
module sky130_sram_4kbyte_1rw_32x1024_8 (
	vccd1,
	vssd1,
	clk0,
	csb0,
	web0,
	wmask0,
	spare_wen0,
	addr0,
	din0,
	dout0
);
	inout vccd1;
	inout vssd1;
	input clk0;
	input csb0;
	input web0;
	input [3:0] wmask0;
	input spare_wen0;
	input [10:0] addr0;
	input [32:0] din0;
	output wire [32:0] dout0;
endmodule
module sky130_sram_0kbytes_1rw_21x64_21 (
	vccd1,
	vssd1,
	clk0,
	csb0,
	web0,
	spare_wen0,
	addr0,
	din0,
	dout0
);
	inout vccd1;
	inout vssd1;
	input clk0;
	input csb0;
	input web0;
	input [6:0] addr0;
	input spare_wen0;
	input [21:0] din0;
	output wire [21:0] dout0;
endmodule